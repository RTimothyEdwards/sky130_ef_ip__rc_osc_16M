VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_ef_ip__rc_osc_16M
  CLASS BLOCK ;
  FOREIGN sky130_ef_ip__rc_osc_16M ;
  ORIGIN 0.000 0.000 ;
  SIZE 61.210 BY 53.620 ;
  PIN avdd
    ANTENNADIFFAREA 137.480896 ;
    PORT
      LAYER met2 ;
        RECT -0.120 38.695 53.690 44.285 ;
    END
    PORT
      LAYER met2 ;
        RECT 54.130 38.695 54.630 44.285 ;
    END
  END avdd
  PIN avss
    ANTENNADIFFAREA 96.482201 ;
    PORT
      LAYER met2 ;
        RECT 52.890 9.720 54.680 15.310 ;
    END
    PORT
      LAYER met2 ;
        RECT -0.120 9.720 1.595 15.310 ;
    END
  END avss
  PIN dvss
    ANTENNADIFFAREA 5.493300 ;
    PORT
      LAYER met1 ;
        RECT 52.540 31.910 54.630 35.795 ;
    END
  END dvss
  PIN dvdd
    ANTENNADIFFAREA 5.371800 ;
    PORT
      LAYER met1 ;
        RECT 52.540 18.170 54.680 23.490 ;
    END
  END dvdd
  PIN ena
    ANTENNAGATEAREA 0.985500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met2 ;
        RECT 53.850 25.070 54.850 26.070 ;
    END
  END ena
  PIN dout
    ANTENNADIFFAREA 0.731800 ;
    PORT
      LAYER met2 ;
        RECT 53.850 29.340 54.850 30.340 ;
    END
  END dout
  OBS
      LAYER nwell ;
        RECT -0.120 3.400 54.885 50.410 ;
      LAYER li1 ;
        RECT 0.310 3.865 54.705 49.970 ;
      LAYER met1 ;
        RECT 0.310 36.075 54.350 47.690 ;
        RECT 0.310 31.630 52.260 36.075 ;
        RECT 0.310 23.770 54.350 31.630 ;
        RECT 0.310 17.890 52.260 23.770 ;
        RECT 0.310 6.090 54.350 17.890 ;
      LAYER met2 ;
        RECT 0.340 44.565 54.285 47.700 ;
        RECT 0.340 30.620 54.285 38.415 ;
        RECT 0.340 29.060 53.570 30.620 ;
        RECT 0.340 26.350 54.285 29.060 ;
        RECT 0.340 24.790 53.570 26.350 ;
        RECT 0.340 15.590 54.285 24.790 ;
        RECT 1.875 9.720 52.610 15.590 ;
  END
END sky130_ef_ip__rc_osc_16M
END LIBRARY

