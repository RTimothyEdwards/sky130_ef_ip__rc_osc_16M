magic
tech sky130A
magscale 1 2
timestamp 1747746856
<< dnwell >>
rect 92 6784 10810 9966
rect 92 3972 8858 6784
rect 92 796 10820 3972
<< nwell >>
rect -24 9760 10926 10082
rect -24 1002 298 9760
rect 10604 6990 10926 9760
rect 5886 6052 6872 6731
rect 8652 6668 10926 6990
rect 5886 5374 6256 6052
rect 8652 4088 8974 6668
rect 10497 4937 10551 5411
rect 8652 3766 10936 4088
rect 10614 1002 10936 3766
rect -24 680 10936 1002
<< nsubdiff >>
rect 10461 5035 10487 5353
<< mvnsubdiff >>
rect 49 9989 10853 10009
rect 49 9955 129 9989
rect 10773 9955 10853 9989
rect 49 9935 10853 9955
rect 49 9929 123 9935
rect 49 833 69 9929
rect 103 833 123 9929
rect 10779 9929 10853 9935
rect 10779 6835 10799 9929
rect 10833 6835 10853 9929
rect 10779 6815 10853 6835
rect 8827 6795 10853 6815
rect 8827 6761 8932 6795
rect 10763 6761 10853 6795
rect 8827 6741 10853 6761
rect 8827 6713 8901 6741
rect 8827 4047 8847 6713
rect 8881 4047 8901 6713
rect 8827 4015 8901 4047
rect 8827 3995 10863 4015
rect 8827 3961 8932 3995
rect 10772 3961 10863 3995
rect 8827 3941 10863 3961
rect 49 827 123 833
rect 10789 3927 10863 3941
rect 10789 833 10809 3927
rect 10843 833 10863 3927
rect 10789 827 10863 833
rect 49 807 10863 827
rect 49 773 129 807
rect 10783 773 10863 807
rect 49 753 10863 773
<< mvnsubdiffcont >>
rect 129 9955 10773 9989
rect 69 833 103 9929
rect 10799 6835 10833 9929
rect 8932 6761 10763 6795
rect 8847 4047 8881 6713
rect 8932 3961 10772 3995
rect 10809 833 10843 3927
rect 129 773 10783 807
<< locali >>
rect 62 9989 10835 9994
rect 62 9955 129 9989
rect 10773 9955 10835 9989
rect 62 9929 10835 9955
rect 62 833 69 9929
rect 103 9851 10799 9929
rect 103 7721 186 9851
rect 169 4023 186 7721
rect 295 9633 10588 9747
rect 295 7128 409 9633
rect 10474 7128 10588 9633
rect 295 7109 10588 7128
rect 295 7024 7186 7109
rect 8627 7024 10588 7109
rect 295 7014 10588 7024
rect 10730 8848 10799 9851
rect 10833 9851 10835 9929
rect 10730 7750 10738 8848
rect 496 7012 1636 7014
rect 496 5331 1174 7012
rect 10730 6911 10799 7750
rect 2181 6769 6769 6770
rect 2134 6743 6769 6769
rect 2134 6686 2219 6743
rect 6746 6686 6769 6743
rect 1294 6611 6769 6686
rect 1294 6168 1448 6611
rect 6449 6169 6769 6611
rect 8739 6884 10799 6911
rect 8739 6859 8915 6884
rect 1852 6168 1903 6169
rect 1294 5942 1903 6168
rect 2177 5942 2503 6168
rect 2777 5942 3119 6168
rect 3393 5942 3735 6168
rect 4009 5942 4351 6168
rect 4625 5942 4967 6168
rect 5241 5942 5583 6168
rect 6449 6168 6893 6169
rect 5857 6095 6893 6168
rect 5857 5942 6349 6095
rect 6760 5942 6893 6095
rect 1294 5487 1448 5942
rect 6765 5487 6893 5942
rect 1294 5330 6893 5487
rect 2181 5329 6893 5330
rect 2181 5328 6784 5329
rect 6761 5224 6884 5225
rect 1020 5065 6884 5224
rect 1020 4629 1151 5065
rect 5475 4636 6337 5065
rect 1020 4467 1122 4629
rect 5475 4625 5680 4636
rect 1278 4623 5680 4625
rect 1278 4466 1661 4623
rect 1916 4466 2217 4623
rect 2472 4466 2773 4623
rect 3028 4466 3329 4623
rect 3584 4466 3885 4623
rect 4140 4466 4441 4623
rect 4696 4466 4997 4623
rect 5252 4467 5680 4623
rect 5836 4625 6337 4636
rect 6761 4625 6884 5065
rect 5836 4467 6884 4625
rect 5252 4466 6884 4467
rect 6761 4031 6884 4466
rect 103 879 186 4023
rect 1131 3981 6884 4031
rect 1131 3946 6789 3981
rect 1131 3891 1183 3946
rect 6742 3891 6789 3946
rect 8739 3961 8764 6859
rect 8829 6819 8915 6859
rect 10141 6835 10799 6884
rect 10141 6819 10833 6835
rect 8829 6795 10833 6819
rect 8829 6761 8932 6795
rect 10763 6761 10833 6795
rect 8829 6749 10833 6761
rect 8829 6713 8888 6749
rect 8829 4047 8847 6713
rect 8881 4047 8888 6713
rect 9403 6591 9808 6598
rect 9403 6462 9517 6591
rect 9403 5960 9808 6462
rect 10480 6268 10933 6270
rect 9077 5752 9808 5960
rect 9336 5539 9808 5752
rect 10475 6267 10933 6268
rect 10475 6140 10507 6267
rect 10711 6140 10933 6267
rect 10475 6137 10933 6140
rect 10475 6041 10618 6137
rect 10475 5978 10500 6041
rect 10607 5978 10618 6041
rect 10475 5815 10618 5978
rect 10475 5740 10933 5815
rect 9072 5495 9808 5539
rect 9072 5252 9387 5495
rect 9723 5494 9808 5495
rect 10421 5660 10933 5701
rect 10421 5406 10521 5660
rect 10628 5658 10933 5660
rect 10421 5210 10485 5406
rect 10421 5073 10521 5210
rect 10421 5072 10622 5073
rect 10421 5069 10937 5072
rect 10421 4996 10938 5069
rect 10460 4994 10938 4996
rect 10141 4844 10461 4975
rect 8829 4035 8888 4047
rect 8829 4010 10843 4035
rect 8829 3995 9014 4010
rect 9822 3995 10843 4010
rect 8829 3961 8932 3995
rect 10772 3961 10843 3995
rect 8739 3934 9014 3961
rect 9822 3934 10843 3961
rect 8739 3927 10843 3934
rect 8739 3911 10809 3927
rect 1131 3872 6789 3891
rect 306 3771 10595 3789
rect 306 3768 5374 3771
rect 306 3689 1862 3768
rect 3521 3692 5374 3768
rect 7033 3692 10595 3771
rect 3521 3689 10595 3692
rect 306 3675 10595 3689
rect 306 3045 420 3675
rect 306 1960 319 3045
rect 413 1960 420 3045
rect 306 1127 420 1960
rect 10481 3046 10595 3675
rect 10481 1961 10484 3046
rect 10578 1961 10595 3046
rect 10481 1127 10595 1961
rect 306 1013 10595 1127
rect 10740 879 10809 3911
rect 103 833 10809 879
rect 62 807 10843 833
rect 62 773 129 807
rect 10783 773 10843 807
<< viali >>
rect 88 4023 103 7721
rect 103 4023 169 7721
rect 7186 7024 8627 7109
rect 10738 7750 10799 8848
rect 10799 7750 10826 8848
rect 2219 6686 6746 6743
rect 7203 6565 8607 6898
rect 1903 5942 2177 6169
rect 2503 5942 2777 6169
rect 3119 5942 3393 6169
rect 3735 5942 4009 6169
rect 4351 5942 4625 6169
rect 4967 5942 5241 6169
rect 5583 5942 5857 6169
rect 1122 4460 1278 4629
rect 1661 4466 1916 4623
rect 2217 4466 2472 4623
rect 2773 4466 3028 4623
rect 3329 4466 3584 4623
rect 3885 4466 4140 4623
rect 4441 4466 4696 4623
rect 4997 4466 5252 4623
rect 5680 4467 5836 4636
rect 1183 3891 6742 3946
rect 7196 3941 8600 4274
rect 8764 3961 8829 6859
rect 8915 6819 10141 6884
rect 9517 6462 9813 6591
rect 10507 6140 10711 6267
rect 10500 5978 10607 6041
rect 10485 5210 10521 5406
rect 9014 3995 9822 4010
rect 9014 3961 9822 3995
rect 9014 3934 9822 3961
rect 1862 3689 3521 3768
rect 5374 3692 7033 3771
rect 319 1960 413 3045
rect 10484 1961 10578 3046
<< metal1 >>
rect 514 9106 750 9538
rect 846 9106 1082 9538
rect 1178 9106 1414 9538
rect 1510 9106 1746 9538
rect 1842 9106 2078 9538
rect 2174 9106 2410 9538
rect 2506 9106 2742 9538
rect 2838 9514 3074 9538
rect 2838 9126 2916 9514
rect 2990 9126 3074 9514
rect 2838 9106 3074 9126
rect 3170 9106 3406 9538
rect 3502 9106 3738 9538
rect 3834 9106 4070 9538
rect 4166 9106 4402 9538
rect 4498 9106 4734 9538
rect 4830 9106 5066 9538
rect 5162 9106 5398 9538
rect 5494 9106 5730 9538
rect 5826 9106 6062 9538
rect 6158 9106 6394 9538
rect 6490 9106 6726 9538
rect 6822 9106 7058 9538
rect 7154 9106 7390 9538
rect 7486 9106 7722 9538
rect 7818 9106 8054 9538
rect 8150 9106 8386 9538
rect 8482 9106 8718 9538
rect 8814 9106 9050 9538
rect 9146 9106 9382 9538
rect 9478 9106 9714 9538
rect 9810 9106 10046 9538
rect 10142 9106 10378 9538
rect 10732 8848 10832 8860
rect 10728 7750 10738 8848
rect 10826 7750 10836 8848
rect 10732 7738 10832 7750
rect 82 7721 175 7733
rect 78 4023 88 7721
rect 169 6481 179 7721
rect 513 6659 588 7639
rect 680 7206 916 7638
rect 1012 7206 1248 7638
rect 1344 7206 1580 7638
rect 1676 7206 1912 7638
rect 2008 7206 2244 7638
rect 2340 7206 2576 7638
rect 2672 7206 2908 7638
rect 3004 7206 3240 7638
rect 3336 7206 3572 7638
rect 3668 7206 3904 7638
rect 4000 7206 4236 7638
rect 4332 7206 4568 7638
rect 4664 7206 4900 7638
rect 4996 7206 5232 7638
rect 5328 7206 5564 7638
rect 5660 7206 5896 7638
rect 5992 7206 6228 7638
rect 6324 7206 6560 7638
rect 6656 7206 6892 7638
rect 6988 7206 7224 7638
rect 7320 7206 7556 7638
rect 7652 7206 7888 7638
rect 7984 7206 8220 7638
rect 8316 7206 8552 7638
rect 8648 7206 8884 7638
rect 8980 7206 9216 7638
rect 9312 7206 9548 7638
rect 9644 7206 9880 7638
rect 9976 7206 10212 7638
rect 627 7118 1828 7121
rect 7169 7118 8652 7128
rect 627 7109 8652 7118
rect 627 7107 7186 7109
rect 627 6980 654 7107
rect 1795 7024 7186 7107
rect 8627 7024 8652 7109
rect 1795 6980 8652 7024
rect 627 6963 8652 6980
rect 807 6962 8652 6963
rect 7169 6939 8652 6962
rect 8721 7037 10178 7062
rect 7169 6898 8651 6939
rect 2137 6836 6797 6866
rect 2137 6771 2190 6836
rect 6770 6771 6797 6836
rect 2137 6743 6797 6771
rect 2137 6686 2219 6743
rect 6746 6686 6797 6743
rect 2137 6676 6797 6686
rect 513 6608 1278 6659
rect 169 5328 1174 6481
rect 169 4023 179 5328
rect 1230 5327 1278 6608
rect 7169 6565 7203 6898
rect 8607 6565 8651 6898
rect 1507 6493 6061 6540
rect 7169 6524 8651 6565
rect 8721 6919 8761 7037
rect 10142 6919 10178 7037
rect 8721 6884 10178 6919
rect 8721 6859 8915 6884
rect 1507 5632 1554 6493
rect 1626 6284 1665 6493
rect 1736 6350 1985 6436
rect 1790 6180 1917 6350
rect 2053 6285 2092 6493
rect 2162 6349 2209 6493
rect 1790 6169 2192 6180
rect 1790 5942 1903 6169
rect 2177 5942 2192 6169
rect 1790 5931 2192 5942
rect 1627 5632 1666 5821
rect 1790 5764 1917 5931
rect 1725 5669 1994 5764
rect 2052 5632 2091 5819
rect 2157 5632 2204 5753
rect 2373 5714 2420 6493
rect 2483 6283 2514 6493
rect 2573 6175 2673 6433
rect 2491 6169 2789 6175
rect 2491 5942 2503 6169
rect 2777 5942 2789 6169
rect 2491 5936 2789 5942
rect 1507 5585 2204 5632
rect 2336 5667 2420 5714
rect 1230 5276 1839 5327
rect 1439 4964 1449 4985
rect 1194 4641 1278 4889
rect 1348 4738 1376 4955
rect 1384 4924 1449 4964
rect 1439 4923 1449 4924
rect 1606 4923 1616 4985
rect 1116 4629 1284 4641
rect 1112 4460 1122 4629
rect 1278 4460 1288 4629
rect 1116 4448 1284 4460
rect 1454 4147 1486 4886
rect 1788 4808 1839 5276
rect 1960 5081 1970 5102
rect 1903 5040 1970 5081
rect 2127 5081 2137 5102
rect 2127 5044 2217 5081
rect 2127 5040 2137 5044
rect 1903 4740 1940 5040
rect 1649 4623 1928 4629
rect 1649 4466 1661 4623
rect 1916 4466 1928 4623
rect 1649 4460 1928 4466
rect 1747 4203 1831 4460
rect 1904 4147 1937 4346
rect 2009 4147 2049 4897
rect 2180 4770 2217 5044
rect 2336 4804 2383 5667
rect 2482 5106 2514 5820
rect 2588 5670 2692 5936
rect 2985 5671 3029 6440
rect 3099 6283 3130 6493
rect 3189 6175 3289 6433
rect 3107 6169 3405 6175
rect 3107 5942 3119 6169
rect 3393 5942 3405 6169
rect 3107 5936 3405 5942
rect 3092 5346 3131 5825
rect 2993 5181 3003 5346
rect 3060 5304 3131 5346
rect 3190 5344 3229 5752
rect 3601 5671 3645 6440
rect 3715 6283 3746 6493
rect 3805 6175 3905 6433
rect 3723 6169 4021 6175
rect 3723 5942 3735 6169
rect 4009 5942 4021 6169
rect 3723 5936 4021 5942
rect 3708 5344 3747 5825
rect 3190 5305 3747 5344
rect 3819 5346 3858 5756
rect 4217 5671 4261 6440
rect 4331 6283 4362 6493
rect 4421 6175 4521 6433
rect 4339 6169 4637 6175
rect 4339 5942 4351 6169
rect 4625 5942 4637 6169
rect 4339 5936 4637 5942
rect 4324 5346 4363 5825
rect 3819 5307 4363 5346
rect 4445 5346 4484 5763
rect 4833 5671 4877 6440
rect 4947 6283 4978 6493
rect 5037 6175 5137 6433
rect 4955 6169 5253 6175
rect 4955 5942 4967 6169
rect 5241 5942 5253 6169
rect 4955 5936 5253 5942
rect 4940 5346 4979 5825
rect 4445 5307 4979 5346
rect 5048 5346 5087 5755
rect 5449 5671 5493 6440
rect 5563 6283 5594 6493
rect 5653 6175 5753 6433
rect 5872 6356 5923 6493
rect 6078 6177 6178 6439
rect 6386 6191 6396 6290
rect 6756 6191 6766 6290
rect 5571 6169 5869 6175
rect 5571 5942 5583 6169
rect 5857 5942 5869 6169
rect 5571 5936 5869 5942
rect 6069 6168 6246 6177
rect 6069 5942 6077 6168
rect 6236 5942 6246 6168
rect 6069 5935 6246 5942
rect 5556 5346 5595 5825
rect 5672 5350 5711 5762
rect 6395 5684 6479 6191
rect 6904 5985 6914 6006
rect 5048 5307 5595 5346
rect 3060 5181 3070 5304
rect 2472 5044 2482 5106
rect 2639 5044 2649 5106
rect 2459 4770 2496 4977
rect 2180 4733 2496 4770
rect 2205 4623 2484 4629
rect 2205 4466 2217 4623
rect 2472 4466 2484 4623
rect 2205 4460 2484 4466
rect 2303 4449 2395 4460
rect 2311 4206 2395 4449
rect 2461 4148 2494 4351
rect 2561 4206 2603 4895
rect 2904 4699 2946 4892
rect 3016 4738 3055 5181
rect 3190 5033 3229 5305
rect 3128 4994 3229 5033
rect 3128 4805 3167 4994
rect 3460 4699 3502 4892
rect 3572 4738 3611 5305
rect 3819 5034 3858 5307
rect 3679 4995 3858 5034
rect 3679 4799 3718 4995
rect 4016 4699 4058 4892
rect 4128 4738 4167 5307
rect 4445 5036 4484 5307
rect 4235 4997 4484 5036
rect 4235 4807 4274 4997
rect 4572 4699 4614 4892
rect 4684 4738 4723 5307
rect 5048 5039 5087 5307
rect 4789 5000 5087 5039
rect 4789 4799 4828 5000
rect 5128 4699 5170 4892
rect 5240 4738 5279 5307
rect 5659 5185 5669 5350
rect 5726 5308 5736 5350
rect 6540 5308 6584 5959
rect 5726 5241 6584 5308
rect 6642 5947 6914 5985
rect 5726 5185 5736 5241
rect 5672 5038 5711 5185
rect 5347 4999 5711 5038
rect 5347 4800 5386 4999
rect 2904 4657 3159 4699
rect 3460 4657 3715 4699
rect 4016 4657 4271 4699
rect 4572 4657 4827 4699
rect 5128 4657 5383 4699
rect 2761 4623 3040 4629
rect 2761 4466 2773 4623
rect 3028 4466 3040 4623
rect 2761 4460 3040 4466
rect 2859 4449 2951 4460
rect 2867 4206 2951 4449
rect 3017 4148 3050 4351
rect 3117 4206 3159 4657
rect 3317 4623 3596 4629
rect 3317 4466 3329 4623
rect 3584 4466 3596 4623
rect 3317 4460 3596 4466
rect 3415 4449 3507 4460
rect 3423 4206 3507 4449
rect 3573 4148 3606 4351
rect 3673 4206 3715 4657
rect 3873 4623 4152 4629
rect 3873 4466 3885 4623
rect 4140 4466 4152 4623
rect 3873 4460 4152 4466
rect 3971 4449 4063 4460
rect 3979 4206 4063 4449
rect 4129 4148 4162 4351
rect 4229 4206 4271 4657
rect 4429 4623 4708 4629
rect 4429 4466 4441 4623
rect 4696 4466 4708 4623
rect 4429 4460 4708 4466
rect 4527 4449 4619 4460
rect 4535 4206 4619 4449
rect 4685 4148 4718 4351
rect 4785 4206 4827 4657
rect 4985 4623 5264 4629
rect 4985 4466 4997 4623
rect 5252 4466 5264 4623
rect 4985 4460 5264 4466
rect 5083 4449 5175 4460
rect 5091 4206 5175 4449
rect 5241 4148 5274 4351
rect 5341 4206 5383 4657
rect 5674 4636 5842 4648
rect 5674 4631 5680 4636
rect 5540 4623 5680 4631
rect 5540 4466 5549 4623
rect 5836 4467 5842 4636
rect 5804 4466 5842 4467
rect 5540 4457 5842 4466
rect 5674 4455 5842 4457
rect 6087 4465 6131 5241
rect 6428 4641 6466 4878
rect 6533 4761 6569 4951
rect 6642 4803 6680 5947
rect 6904 5928 6914 5947
rect 7105 5928 7115 6006
rect 6934 5163 7307 5197
rect 6934 4979 6968 5163
rect 6814 4915 6824 4979
rect 7011 4915 7021 4979
rect 6533 4725 6956 4761
rect 6917 4656 6956 4725
rect 6428 4603 6679 4641
rect 6917 4617 6981 4656
rect 5708 4292 5792 4455
rect 6087 4422 6574 4465
rect 6218 4421 6574 4422
rect 5708 4291 6468 4292
rect 5708 4209 6478 4291
rect 5708 4208 6366 4209
rect 1454 4099 5518 4147
rect 6530 4142 6574 4421
rect 6641 4208 6679 4603
rect 6971 4592 6981 4617
rect 7168 4592 7178 4656
rect 8721 4334 8764 6859
rect 8609 4324 8764 4334
rect 7152 4274 8764 4324
rect 82 4011 175 4023
rect 1129 3946 6787 4031
rect 1129 3891 1183 3946
rect 6742 3891 6787 3946
rect 7152 3941 7196 4274
rect 8600 3961 8764 4274
rect 8829 6819 8915 6859
rect 10141 6819 10178 6884
rect 8829 6792 10178 6819
rect 8829 4036 8898 6792
rect 10302 6720 10377 7645
rect 9378 6645 10377 6720
rect 9151 6501 9161 6573
rect 9337 6501 9347 6573
rect 9138 6006 9191 6206
rect 9275 6120 9337 6501
rect 8949 5934 8959 6006
rect 9135 5952 9191 6006
rect 9135 5934 9145 5952
rect 9236 5798 9268 6082
rect 9124 5726 9134 5798
rect 9310 5726 9320 5798
rect 9236 5659 9268 5661
rect 9096 5587 9106 5659
rect 9282 5587 9292 5659
rect 9378 4149 9453 6645
rect 9505 6591 9825 6597
rect 9505 6462 9517 6591
rect 9813 6462 9825 6591
rect 10508 6582 10926 7159
rect 9505 6456 9825 6462
rect 10026 6572 10926 6582
rect 10026 6473 10037 6572
rect 10397 6473 10926 6572
rect 10026 6382 10926 6473
rect 9522 6195 9532 6294
rect 9892 6195 9902 6294
rect 10026 6267 10723 6382
rect 9528 4952 9690 6195
rect 10026 6140 10507 6267
rect 10711 6140 10723 6267
rect 10026 6134 10723 6140
rect 10026 6057 10615 6134
rect 10026 6041 10722 6057
rect 10026 5978 10500 6041
rect 10607 5978 10722 6041
rect 10822 6007 10870 6062
rect 10026 5963 10722 5978
rect 10026 5961 10226 5963
rect 10713 5962 10722 5963
rect 10702 5847 10788 5901
rect 10702 5690 10743 5847
rect 10820 5800 10870 6007
rect 10373 5673 10383 5690
rect 10312 5618 10383 5673
rect 10559 5632 10743 5690
rect 10559 5618 10569 5632
rect 10312 5308 10350 5618
rect 10633 5599 10699 5632
rect 10771 5631 10781 5800
rect 10850 5640 10870 5800
rect 10850 5631 10860 5640
rect 10479 5406 10599 5418
rect 10222 5270 10350 5308
rect 10222 5154 10260 5270
rect 10387 5240 10485 5406
rect 10319 5210 10485 5240
rect 10521 5210 10599 5406
rect 10819 5229 10860 5631
rect 10319 5158 10599 5210
rect 10137 5044 10147 5116
rect 10323 5044 10333 5116
rect 10387 4952 10599 5158
rect 10744 4968 10780 5153
rect 9528 4752 10599 4952
rect 10661 4909 10671 4968
rect 10857 4909 10867 4968
rect 10039 4698 10599 4752
rect 10039 4209 10936 4698
rect 9378 4074 10397 4149
rect 8829 4010 9900 4036
rect 8829 3961 9014 4010
rect 8600 3941 9014 3961
rect 7152 3934 9014 3941
rect 9822 3934 9900 4010
rect 7152 3910 9900 3934
rect 1129 3874 6787 3891
rect 1850 3768 3533 3774
rect 1850 3689 1862 3768
rect 3521 3689 3533 3768
rect 1850 3683 3533 3689
rect 5362 3771 7045 3777
rect 5362 3692 5374 3771
rect 7033 3692 7045 3771
rect 5362 3686 7045 3692
rect 62 3543 605 3550
rect 62 3134 76 3543
rect 351 3134 605 3543
rect 62 3118 605 3134
rect 700 3118 936 3550
rect 1032 3118 1268 3550
rect 1364 3118 1600 3550
rect 1696 3118 1932 3550
rect 2028 3118 2264 3550
rect 2360 3118 2596 3550
rect 2692 3118 2928 3550
rect 3024 3118 3260 3550
rect 3356 3118 3592 3550
rect 3688 3118 3924 3550
rect 4020 3118 4256 3550
rect 4352 3118 4588 3550
rect 4684 3118 4920 3550
rect 5016 3118 5252 3550
rect 5348 3118 5584 3550
rect 5680 3118 5916 3550
rect 6012 3118 6248 3550
rect 6344 3118 6580 3550
rect 6676 3118 6912 3550
rect 7008 3118 7244 3550
rect 7340 3118 7576 3550
rect 7672 3118 7908 3550
rect 8004 3118 8240 3550
rect 8336 3118 8572 3550
rect 8668 3118 8904 3550
rect 9000 3118 9236 3550
rect 9332 3118 9568 3550
rect 9664 3118 9900 3550
rect 9996 3118 10232 3550
rect 10322 3115 10397 4074
rect 10508 3634 10936 4209
rect 313 3045 419 3057
rect 10478 3046 10584 3058
rect 309 1960 319 3045
rect 413 1960 423 3045
rect 10474 1961 10484 3046
rect 10578 1961 10588 3046
rect 313 1948 419 1960
rect 10478 1949 10584 1961
rect 534 1218 770 1650
rect 866 1218 1102 1650
rect 1198 1218 1434 1650
rect 1530 1218 1766 1650
rect 1862 1218 2098 1650
rect 2194 1218 2430 1650
rect 2526 1218 2762 1650
rect 2858 1218 3094 1650
rect 3190 1218 3426 1650
rect 3522 1218 3758 1650
rect 3854 1218 4090 1650
rect 4186 1218 4422 1650
rect 4518 1218 4754 1650
rect 4850 1218 5086 1650
rect 5182 1218 5418 1650
rect 5514 1218 5750 1650
rect 5846 1218 6082 1650
rect 6178 1218 6414 1650
rect 6510 1218 6746 1650
rect 6842 1218 7078 1650
rect 7174 1218 7410 1650
rect 7506 1218 7742 1650
rect 7838 1218 8074 1650
rect 8170 1218 8406 1650
rect 8502 1218 8738 1650
rect 8834 1218 9070 1650
rect 9166 1218 9402 1650
rect 9498 1218 9734 1650
rect 9830 1218 10066 1650
rect 10162 1218 10398 1650
<< via1 >>
rect 2916 9126 2990 9514
rect 10738 7750 10826 8848
rect 88 4023 169 7721
rect 654 6980 1795 7107
rect 2190 6771 6770 6836
rect 7203 6565 8607 6898
rect 8761 6919 10142 7037
rect 2503 5942 2777 6169
rect 1449 4923 1606 4985
rect 1122 4460 1278 4629
rect 1970 5040 2127 5102
rect 1661 4466 1916 4623
rect 3119 5942 3393 6169
rect 3003 5181 3060 5346
rect 3735 5942 4009 6169
rect 4351 5942 4625 6169
rect 4967 5942 5241 6169
rect 6396 6191 6756 6290
rect 5583 5942 5857 6169
rect 6077 5942 6236 6168
rect 2482 5044 2639 5106
rect 2217 4466 2472 4623
rect 5669 5185 5726 5350
rect 2773 4466 3028 4623
rect 3329 4466 3584 4623
rect 3885 4466 4140 4623
rect 4441 4466 4696 4623
rect 4997 4466 5252 4623
rect 5549 4467 5680 4623
rect 5680 4467 5804 4623
rect 5549 4466 5804 4467
rect 6914 5928 7105 6006
rect 6824 4915 7011 4979
rect 6981 4592 7168 4656
rect 1183 3891 6742 3946
rect 7196 3941 8600 4274
rect 9161 6501 9337 6573
rect 8959 5934 9135 6006
rect 9134 5726 9310 5798
rect 9106 5587 9282 5659
rect 9517 6462 9813 6591
rect 10037 6473 10397 6572
rect 9532 6195 9892 6294
rect 10383 5618 10559 5690
rect 10781 5631 10850 5800
rect 9871 5040 9930 5226
rect 10147 5044 10323 5116
rect 10671 4909 10857 4968
rect 1862 3689 3521 3768
rect 5374 3692 7033 3771
rect 76 3134 351 3543
rect 319 1960 413 3045
rect 10484 1961 10578 3046
<< metal2 >>
rect 2838 9514 3074 9540
rect 2838 9126 2916 9514
rect 2990 9126 3074 9514
rect 2838 8857 3074 9126
rect 10738 8857 10826 8858
rect -24 8848 10926 8857
rect -24 7750 10738 8848
rect 10826 7750 10926 8848
rect -24 7739 10926 7750
rect 68 7721 358 7739
rect 68 4023 88 7721
rect 169 4023 358 7721
rect 627 7107 1828 7121
rect 627 7103 654 7107
rect 68 3543 358 4023
rect 68 3134 76 3543
rect 351 3134 358 3543
rect 68 3128 358 3134
rect 625 6980 654 7103
rect 1795 6980 1828 7107
rect 625 6963 1828 6980
rect 625 6896 1175 6963
rect 625 5312 1174 6896
rect 2453 6883 4111 7739
rect 5409 6889 5980 7739
rect 9837 7194 10178 7739
rect 7169 6939 8652 7128
rect 8721 7037 10178 7194
rect 7169 6898 8651 6939
rect 8721 6919 8761 7037
rect 10142 6919 10178 7037
rect 8721 6900 10178 6919
rect 5409 6883 6838 6889
rect 2119 6836 6838 6883
rect 2119 6771 2190 6836
rect 6770 6771 6838 6836
rect 2119 6673 6838 6771
rect 2453 6217 4111 6673
rect 5409 6217 5951 6673
rect 7169 6565 7203 6898
rect 8607 6565 8651 6898
rect 9517 6592 9813 6601
rect 7169 6524 8651 6565
rect 9147 6591 10402 6592
rect 9147 6573 9517 6591
rect 9147 6501 9161 6573
rect 9337 6501 9517 6573
rect 9147 6462 9517 6501
rect 9813 6572 10402 6591
rect 9813 6473 10037 6572
rect 10397 6473 10402 6572
rect 9813 6462 10402 6473
rect 9147 6460 10402 6462
rect 9517 6452 9813 6460
rect 6396 6292 6756 6300
rect 9532 6294 9892 6304
rect 6396 6290 9532 6292
rect 1538 6169 6284 6217
rect 6756 6195 9532 6290
rect 6756 6194 9892 6195
rect 6396 6181 6756 6191
rect 9532 6185 9892 6194
rect 1538 5942 2503 6169
rect 2777 5942 3119 6169
rect 3393 5942 3735 6169
rect 4009 5942 4351 6169
rect 4625 5942 4967 6169
rect 5241 5942 5583 6169
rect 5857 6168 6284 6169
rect 5857 5942 6077 6168
rect 6236 5942 6284 6168
rect 1538 5901 6284 5942
rect 6914 6006 7105 6016
rect 8959 6006 9135 6016
rect 7105 5947 8856 5991
rect 8958 5947 8959 5991
rect 6914 5918 7105 5928
rect 8812 5894 8856 5947
rect 10770 5991 10970 6068
rect 9135 5947 10970 5991
rect 8959 5924 9135 5934
rect 8812 5850 10308 5894
rect 10770 5868 10970 5947
rect 9134 5798 9310 5808
rect 9134 5716 9310 5726
rect 10264 5672 10308 5850
rect 10781 5800 10850 5868
rect 10383 5690 10559 5700
rect 9106 5659 9282 5669
rect 3003 5346 3060 5356
rect 625 4662 1175 5312
rect 5669 5350 5726 5360
rect 3060 5238 5669 5279
rect 3003 5171 3060 5181
rect 5669 5175 5726 5185
rect 1970 5102 2127 5112
rect 2482 5106 2639 5116
rect 1932 5041 1970 5102
rect 2127 5044 2482 5102
rect 2639 5044 7147 5102
rect 2127 5041 7147 5044
rect 1970 5030 2127 5040
rect 2482 5034 2639 5041
rect 1449 4985 1606 4995
rect 6814 4979 7011 4989
rect 6814 4968 6824 4979
rect 1606 4923 6824 4968
rect 1449 4913 1606 4923
rect 6824 4905 7011 4915
rect 7086 4944 7147 5041
rect 7086 4883 7916 4944
rect 625 4629 6019 4662
rect 6981 4657 7168 4666
rect 8572 4657 8637 5618
rect 10264 5628 10383 5672
rect 10781 5621 10850 5631
rect 10383 5608 10559 5618
rect 9106 5577 9282 5587
rect 9900 5409 10453 5463
rect 9863 5040 9871 5226
rect 9930 5040 9939 5226
rect 10147 5116 10323 5126
rect 10399 5104 10453 5409
rect 10323 5071 10453 5104
rect 10770 5071 10970 5214
rect 10323 5057 10970 5071
rect 9871 4969 9930 5040
rect 10147 5034 10323 5044
rect 10399 5017 10970 5057
rect 10770 5014 10970 5017
rect 10671 4969 10857 4976
rect 9871 4968 10857 4969
rect 9871 4910 10671 4968
rect 10671 4899 10857 4909
rect 625 4460 1122 4629
rect 1278 4623 6019 4629
rect 1278 4466 1661 4623
rect 1916 4466 2217 4623
rect 2472 4466 2773 4623
rect 3028 4466 3329 4623
rect 3584 4466 3885 4623
rect 4140 4466 4441 4623
rect 4696 4466 4997 4623
rect 5252 4466 5549 4623
rect 5804 4466 6019 4623
rect 6979 4656 8637 4657
rect 6979 4592 6981 4656
rect 7168 4592 8637 4656
rect 6981 4582 7168 4592
rect 1278 4460 6019 4466
rect 625 4360 6019 4460
rect 625 4056 1175 4360
rect 1861 4056 3520 4360
rect 5375 4056 5918 4360
rect 7152 4274 8634 4324
rect 625 3946 6814 4056
rect 625 3891 1183 3946
rect 6742 3891 6814 3946
rect 7152 3941 7196 4274
rect 8600 3941 8634 4274
rect 7152 3910 8634 3941
rect 625 3842 6814 3891
rect 625 3062 1175 3842
rect 1861 3768 3521 3842
rect 1861 3689 1862 3768
rect 1861 3679 3521 3689
rect 5374 3771 7034 3842
rect 7033 3692 7034 3771
rect 5374 3682 7034 3692
rect 1861 3062 3520 3679
rect 5375 3654 7034 3682
rect 5375 3062 5905 3654
rect 6213 3062 6971 3654
rect -24 3046 10936 3062
rect -24 3045 10484 3046
rect -24 1960 319 3045
rect 413 1961 10484 3045
rect 10578 1961 10936 3046
rect 413 1960 10936 1961
rect -24 1944 10936 1960
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D3 paramcells
timestamp 1699295625
transform 1 0 9223 0 1 5622
box -183 -183 183 183
use rc_osc_level_shifter  rc_osc_level_shifter_0
timestamp 1699295625
transform -1 0 9816 0 -1 4232
box -422 -2544 2736 144
use sky130_fd_pr__nfet_01v8_L9WNCD  sky130_fd_pr__nfet_01v8_L9WNCD_0 paramcells
timestamp 1699295625
transform 1 0 10759 0 1 5976
box -211 -229 211 229
use sky130_fd_pr__pfet_01v8_2Z69BZ  sky130_fd_pr__pfet_01v8_2Z69BZ_0 paramcells
timestamp 1699295625
transform 1 0 10286 0 1 5163
box -211 -226 211 226
use sky130_fd_pr__pfet_01v8_856REK  sky130_fd_pr__pfet_01v8_856REK_0 paramcells
timestamp 1716055179
transform 1 0 10714 0 -1 5368
box -263 -369 263 369
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  sky130_fd_pr__pfet_g5v0d10v5_6ELFTH_0 paramcells
timestamp 1699295625
transform 1 0 2498 0 1 6391
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  sky130_fd_pr__pfet_g5v0d10v5_6ELFTH_1
timestamp 1699295625
transform 1 0 1646 0 1 6391
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  sky130_fd_pr__pfet_g5v0d10v5_6ELFTH_2
timestamp 1699295625
transform 1 0 2072 0 1 6391
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  sky130_fd_pr__pfet_g5v0d10v5_6ELFTH_3
timestamp 1699295625
transform 1 0 2498 0 1 5713
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  sky130_fd_pr__pfet_g5v0d10v5_6ELFTH_4
timestamp 1699295625
transform 1 0 2072 0 1 5713
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  sky130_fd_pr__pfet_g5v0d10v5_6ELFTH_5
timestamp 1699295625
transform 1 0 5578 0 1 6391
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_T537S5  sky130_fd_pr__pfet_g5v0d10v5_T537S5_0 paramcells
timestamp 1716055179
transform 1 0 6560 0 1 5770
box -308 -423 308 423
use sky130_fd_pr__res_xhigh_po_0p35_NVJ5PF  sky130_fd_pr__res_xhigh_po_0p35_NVJ5PF_0 paramcells
timestamp 1715996061
transform 1 0 5466 0 1 2384
box -5098 -1332 5098 1332
use sky130_fd_pr__res_xhigh_po_0p35_NVJ5PF  sky130_fd_pr__res_xhigh_po_0p35_NVJ5PF_1
timestamp 1715996061
transform 1 0 5446 0 1 8372
box -5098 -1332 5098 1332
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM1 paramcells
timestamp 1699295625
transform 1 0 3032 0 1 4848
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM2
timestamp 1699295625
transform 1 0 3114 0 1 5713
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM3
timestamp 1699295625
transform 1 0 3730 0 1 5713
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM4
timestamp 1699295625
transform 1 0 3588 0 1 4848
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM7
timestamp 1699295625
transform 1 0 4962 0 1 5713
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM8
timestamp 1699295625
transform 1 0 4700 0 1 4848
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM9
timestamp 1699295625
transform 1 0 4346 0 1 5713
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM10
timestamp 1699295625
transform 1 0 4144 0 1 4848
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM12
timestamp 1699295625
transform 1 0 6552 0 1 4246
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM13
timestamp 1699295625
transform 1 0 6552 0 1 4846
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM15
timestamp 1699295625
transform 1 0 5578 0 1 5713
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM16
timestamp 1699295625
transform 1 0 5256 0 1 4848
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM17
timestamp 1699295625
transform 1 0 4962 0 1 6391
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM18
timestamp 1699295625
transform 1 0 6004 0 1 6391
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM19
timestamp 1699295625
transform 1 0 5256 0 1 4248
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM20
timestamp 1699295625
transform 1 0 4700 0 1 4248
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM21
timestamp 1699295625
transform 1 0 1920 0 1 4248
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM23
timestamp 1699295625
transform 1 0 1920 0 1 4846
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM24
timestamp 1699295625
transform 1 0 3114 0 1 6391
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM25
timestamp 1699295625
transform 1 0 3730 0 1 6391
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM26
timestamp 1699295625
transform 1 0 4346 0 1 6391
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM27
timestamp 1699295625
transform 1 0 4144 0 1 4248
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM28
timestamp 1699295625
transform 1 0 3588 0 1 4248
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM29
timestamp 1699295625
transform 1 0 3032 0 1 4248
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM30
timestamp 1699295625
transform 1 0 2476 0 1 4248
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM33
timestamp 1699295625
transform 1 0 1364 0 1 4846
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM34
timestamp 1699295625
transform 1 0 1646 0 1 5713
box -308 -339 308 339
use sky130_fd_pr__nfet_01v8_L7BSKG  XM35 paramcells
timestamp 1699295625
transform 1 0 9251 0 1 6131
box -211 -221 211 221
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM36
timestamp 1699295625
transform 1 0 2476 0 1 4848
box -278 -300 278 300
<< labels >>
flabel metal2 s 10578 1944 10886 3062 0 FreeSans 960 90 0 0 avss
port 1 nsew
flabel metal1 10736 3634 10936 4391 0 FreeSans 256 0 0 0 dvdd
port 3 nsew
flabel metal2 -24 1944 176 3062 0 FreeSans 256 0 0 0 avss
port 1 nsew
flabel metal1 10726 6382 10926 7139 0 FreeSans 256 0 0 0 dvss
port 2 nsew
flabel metal2 10770 5014 10970 5214 0 FreeSans 256 0 0 0 ena
port 4 nsew
flabel metal2 10770 5868 10970 6068 0 FreeSans 256 0 0 0 dout
port 5 nsew
flabel metal2 -24 7739 176 8857 0 FreeSans 256 0 0 0 avdd
port 0 nsew
flabel metal2 s 10826 7739 10926 8857 0 FreeSans 640 90 0 0 avdd
port 0 nsew
<< properties >>
string FIXED_BBOX 0 0 12242 10724
<< end >>
