magic
tech sky130A
magscale 1 2
timestamp 1716066989
<< dnwell >>
rect 116 6766 10770 9908
rect 116 3954 8858 6766
rect 116 816 10770 3954
<< nwell >>
rect 0 9702 10886 10024
rect 0 1022 322 9702
rect 10564 6972 10886 9702
rect 5886 6034 6872 6713
rect 8652 6650 10886 6972
rect 5886 5356 6256 6034
rect 8652 4070 8974 6650
rect 10497 4919 10551 5393
rect 8652 3805 10886 4070
rect 9768 3748 10886 3805
rect 10564 1022 10886 3748
rect 0 700 10886 1022
<< nsubdiff >>
rect 10461 5017 10487 5335
<< mvnsubdiff >>
rect 73 9931 10813 9951
rect 73 9897 153 9931
rect 10733 9897 10813 9931
rect 73 9877 10813 9897
rect 73 9871 147 9877
rect 73 853 93 9871
rect 127 853 147 9871
rect 10739 9871 10813 9877
rect 10739 6817 10759 9871
rect 10793 6817 10813 9871
rect 10739 6797 10813 6817
rect 8827 6777 10813 6797
rect 8827 6743 8932 6777
rect 10723 6743 10813 6777
rect 8827 6723 10813 6743
rect 8827 6695 8901 6723
rect 8827 4029 8847 6695
rect 8881 4029 8901 6695
rect 8827 3997 8901 4029
rect 8827 3977 10813 3997
rect 8827 3943 8932 3977
rect 10722 3943 10813 3977
rect 8827 3923 10813 3943
rect 73 847 147 853
rect 10739 3909 10813 3923
rect 10739 853 10759 3909
rect 10793 853 10813 3909
rect 10739 847 10813 853
rect 73 827 10813 847
rect 73 793 153 827
rect 10733 793 10813 827
rect 73 773 10813 793
<< mvnsubdiffcont >>
rect 153 9897 10733 9931
rect 93 853 127 9871
rect 10759 6817 10793 9871
rect 8932 6743 10723 6777
rect 8847 4029 8881 6695
rect 8932 3943 10722 3977
rect 10759 853 10793 3909
rect 153 793 10733 827
<< locali >>
rect 86 9931 10795 9936
rect 86 9897 153 9931
rect 10733 9897 10795 9931
rect 86 9871 10795 9897
rect 86 853 93 9871
rect 127 9793 10759 9871
rect 127 7683 210 9793
rect 193 4005 210 7683
rect 295 9595 10588 9709
rect 295 7090 409 9595
rect 10474 7090 10588 9595
rect 295 7071 10588 7090
rect 295 6986 7186 7071
rect 8627 6986 10588 7071
rect 295 6976 10588 6986
rect 10690 8810 10759 9793
rect 10793 9793 10795 9871
rect 10690 7712 10698 8810
rect 496 6974 1636 6976
rect 496 5313 1174 6974
rect 10690 6893 10759 7712
rect 2181 6751 6769 6752
rect 2134 6725 6769 6751
rect 2134 6668 2219 6725
rect 6746 6668 6769 6725
rect 1294 6593 6769 6668
rect 1294 6150 1448 6593
rect 6449 6151 6769 6593
rect 8739 6866 10759 6893
rect 8739 6841 8915 6866
rect 1852 6150 1903 6151
rect 1294 5924 1903 6150
rect 2177 5924 2503 6150
rect 2777 5924 3119 6150
rect 3393 5924 3735 6150
rect 4009 5924 4351 6150
rect 4625 5924 4967 6150
rect 5241 5924 5583 6150
rect 6449 6150 6893 6151
rect 5857 6077 6893 6150
rect 5857 5924 6349 6077
rect 6760 5924 6893 6077
rect 1294 5469 1448 5924
rect 6765 5469 6893 5924
rect 1294 5312 6893 5469
rect 2181 5311 6893 5312
rect 2181 5310 6784 5311
rect 6761 5206 6884 5207
rect 1020 5047 6884 5206
rect 1020 4611 1151 5047
rect 5475 4618 6337 5047
rect 1020 4449 1122 4611
rect 5475 4607 5680 4618
rect 1278 4605 5680 4607
rect 1278 4448 1661 4605
rect 1916 4448 2217 4605
rect 2472 4448 2773 4605
rect 3028 4448 3329 4605
rect 3584 4448 3885 4605
rect 4140 4448 4441 4605
rect 4696 4448 4997 4605
rect 5252 4449 5680 4605
rect 5836 4607 6337 4618
rect 6761 4607 6884 5047
rect 5836 4449 6884 4607
rect 5252 4448 6884 4449
rect 6761 4013 6884 4448
rect 127 899 210 4005
rect 1131 3963 6884 4013
rect 1131 3928 6789 3963
rect 1131 3873 1183 3928
rect 6742 3873 6789 3928
rect 8739 3943 8764 6841
rect 8829 6801 8915 6841
rect 10141 6817 10759 6866
rect 10141 6801 10793 6817
rect 8829 6777 10793 6801
rect 8829 6743 8932 6777
rect 10723 6743 10793 6777
rect 8829 6731 10793 6743
rect 8829 6695 8888 6731
rect 8829 4029 8847 6695
rect 8881 4029 8888 6695
rect 9403 6573 9808 6580
rect 9403 6444 9517 6573
rect 9403 5942 9808 6444
rect 10480 6250 10933 6252
rect 9077 5734 9808 5942
rect 9336 5521 9808 5734
rect 10475 6249 10933 6250
rect 10475 6122 10507 6249
rect 10711 6122 10933 6249
rect 10475 6119 10933 6122
rect 10475 6023 10618 6119
rect 10475 5960 10500 6023
rect 10607 5960 10618 6023
rect 10475 5797 10618 5960
rect 10475 5722 10933 5797
rect 9072 5477 9808 5521
rect 9072 5234 9387 5477
rect 9723 5476 9808 5477
rect 10421 5642 10933 5683
rect 10421 5388 10521 5642
rect 10628 5640 10933 5642
rect 10421 5192 10485 5388
rect 10421 5055 10521 5192
rect 10421 5054 10622 5055
rect 10421 5051 10937 5054
rect 10421 4978 10938 5051
rect 10460 4976 10938 4978
rect 10141 4826 10461 4957
rect 8829 4017 8888 4029
rect 8829 3977 10793 4017
rect 8829 3943 8932 3977
rect 10722 3943 10793 3977
rect 8739 3909 10793 3943
rect 8739 3893 10759 3909
rect 1131 3854 6789 3873
rect 306 3771 10595 3789
rect 306 3768 5374 3771
rect 306 3689 1862 3768
rect 3521 3692 5374 3768
rect 7033 3692 10595 3771
rect 3521 3689 10595 3692
rect 306 3675 10595 3689
rect 306 3045 420 3675
rect 306 1960 319 3045
rect 413 1960 420 3045
rect 306 1127 420 1960
rect 10481 3046 10595 3675
rect 10481 1961 10484 3046
rect 10578 1961 10595 3046
rect 10481 1127 10595 1961
rect 306 1013 10595 1127
rect 10690 899 10759 3893
rect 127 853 10759 899
rect 86 827 10793 853
rect 86 793 153 827
rect 10733 793 10793 827
<< viali >>
rect 112 4005 127 7683
rect 127 4005 193 7683
rect 7186 6986 8627 7071
rect 10698 7712 10759 8810
rect 10759 7712 10786 8810
rect 2219 6668 6746 6725
rect 7203 6547 8607 6880
rect 1903 5924 2177 6151
rect 2503 5924 2777 6151
rect 3119 5924 3393 6151
rect 3735 5924 4009 6151
rect 4351 5924 4625 6151
rect 4967 5924 5241 6151
rect 5583 5924 5857 6151
rect 1122 4442 1278 4611
rect 1661 4448 1916 4605
rect 2217 4448 2472 4605
rect 2773 4448 3028 4605
rect 3329 4448 3584 4605
rect 3885 4448 4140 4605
rect 4441 4448 4696 4605
rect 4997 4448 5252 4605
rect 5680 4449 5836 4618
rect 1183 3873 6742 3928
rect 7196 3923 8600 4256
rect 8764 3943 8829 6841
rect 8915 6801 10141 6866
rect 9517 6444 9813 6573
rect 10507 6122 10711 6249
rect 10500 5960 10607 6023
rect 10485 5192 10521 5388
rect 1862 3689 3521 3768
rect 5374 3692 7033 3771
rect 319 1960 413 3045
rect 10484 1961 10578 3046
<< metal1 >>
rect 514 9068 750 9500
rect 846 9068 1082 9500
rect 1178 9068 1414 9500
rect 1510 9068 1746 9500
rect 1842 9068 2078 9500
rect 2174 9068 2410 9500
rect 2506 9068 2742 9500
rect 2838 9068 3074 9500
rect 3170 9068 3406 9500
rect 3502 9068 3738 9500
rect 3834 9068 4070 9500
rect 4166 9068 4402 9500
rect 4498 9068 4734 9500
rect 4830 9068 5066 9500
rect 5162 9068 5398 9500
rect 5494 9068 5730 9500
rect 5826 9068 6062 9500
rect 6158 9068 6394 9500
rect 6490 9068 6726 9500
rect 6822 9068 7058 9500
rect 7154 9068 7390 9500
rect 7486 9068 7722 9500
rect 7818 9068 8054 9500
rect 8150 9068 8386 9500
rect 8482 9068 8718 9500
rect 8814 9068 9050 9500
rect 9146 9068 9382 9500
rect 9478 9068 9714 9500
rect 9810 9068 10046 9500
rect 10142 9068 10378 9500
rect 10692 8810 10792 8822
rect 10688 7712 10698 8810
rect 10786 7712 10796 8810
rect 10692 7700 10792 7712
rect 106 7683 199 7695
rect 102 4005 112 7683
rect 193 6463 203 7683
rect 513 6641 588 7601
rect 680 7168 916 7600
rect 1012 7168 1248 7600
rect 1344 7168 1580 7600
rect 1676 7168 1912 7600
rect 2008 7168 2244 7600
rect 2340 7168 2576 7600
rect 2672 7168 2908 7600
rect 3004 7168 3240 7600
rect 3336 7168 3572 7600
rect 3668 7168 3904 7600
rect 4000 7168 4236 7600
rect 4332 7168 4568 7600
rect 4664 7168 4900 7600
rect 4996 7168 5232 7600
rect 5328 7168 5564 7600
rect 5660 7168 5896 7600
rect 5992 7168 6228 7600
rect 6324 7168 6560 7600
rect 6656 7168 6892 7600
rect 6988 7168 7224 7600
rect 7320 7168 7556 7600
rect 7652 7168 7888 7600
rect 7984 7168 8220 7600
rect 8316 7168 8552 7600
rect 8648 7168 8884 7600
rect 8980 7168 9216 7600
rect 9312 7168 9548 7600
rect 9644 7168 9880 7600
rect 9976 7168 10212 7600
rect 627 7080 1828 7083
rect 7169 7080 8652 7090
rect 627 7071 8652 7080
rect 627 7069 7186 7071
rect 627 6942 654 7069
rect 1795 6986 7186 7069
rect 8627 6986 8652 7071
rect 1795 6942 8652 6986
rect 627 6925 8652 6942
rect 807 6924 8652 6925
rect 7169 6901 8652 6924
rect 8721 6999 10178 7024
rect 8721 6901 8761 6999
rect 10142 6901 10178 6999
rect 7169 6880 8651 6901
rect 2137 6818 6797 6848
rect 2137 6753 2190 6818
rect 6770 6753 6797 6818
rect 2137 6725 6797 6753
rect 2137 6668 2219 6725
rect 6746 6668 6797 6725
rect 2137 6658 6797 6668
rect 513 6590 1278 6641
rect 193 5310 1174 6463
rect 193 4005 203 5310
rect 1230 5309 1278 6590
rect 7169 6547 7203 6880
rect 8607 6547 8651 6880
rect 1507 6475 6061 6522
rect 7169 6506 8651 6547
rect 8721 6866 10178 6901
rect 8721 6841 8915 6866
rect 1507 5614 1554 6475
rect 1626 6266 1665 6475
rect 1736 6332 1985 6418
rect 1790 6162 1917 6332
rect 2053 6267 2092 6475
rect 2162 6331 2209 6475
rect 1790 6151 2192 6162
rect 1790 5924 1903 6151
rect 2177 5924 2192 6151
rect 1790 5913 2192 5924
rect 1627 5614 1666 5803
rect 1790 5746 1917 5913
rect 1725 5651 1994 5746
rect 2052 5614 2091 5801
rect 2157 5614 2204 5735
rect 2373 5696 2420 6475
rect 2483 6265 2514 6475
rect 2573 6157 2673 6415
rect 2491 6151 2789 6157
rect 2491 5924 2503 6151
rect 2777 5924 2789 6151
rect 2491 5918 2789 5924
rect 1507 5567 2204 5614
rect 2336 5649 2420 5696
rect 1230 5258 1839 5309
rect 1439 4946 1449 4967
rect 1194 4623 1278 4871
rect 1348 4720 1376 4937
rect 1384 4906 1449 4946
rect 1439 4905 1449 4906
rect 1606 4905 1616 4967
rect 1116 4611 1284 4623
rect 1112 4442 1122 4611
rect 1278 4442 1288 4611
rect 1116 4430 1284 4442
rect 1454 4129 1486 4868
rect 1788 4790 1839 5258
rect 1960 5063 1970 5084
rect 1903 5022 1970 5063
rect 2127 5063 2137 5084
rect 2127 5026 2217 5063
rect 2127 5022 2137 5026
rect 1903 4722 1940 5022
rect 1649 4605 1928 4611
rect 1649 4448 1661 4605
rect 1916 4448 1928 4605
rect 1649 4442 1928 4448
rect 1747 4185 1831 4442
rect 1904 4129 1937 4328
rect 2009 4129 2049 4879
rect 2180 4752 2217 5026
rect 2336 4786 2383 5649
rect 2482 5088 2514 5802
rect 2588 5652 2692 5918
rect 2985 5653 3029 6422
rect 3099 6265 3130 6475
rect 3189 6157 3289 6415
rect 3107 6151 3405 6157
rect 3107 5924 3119 6151
rect 3393 5924 3405 6151
rect 3107 5918 3405 5924
rect 3092 5328 3131 5807
rect 2993 5163 3003 5328
rect 3060 5286 3131 5328
rect 3190 5326 3229 5734
rect 3601 5653 3645 6422
rect 3715 6265 3746 6475
rect 3805 6157 3905 6415
rect 3723 6151 4021 6157
rect 3723 5924 3735 6151
rect 4009 5924 4021 6151
rect 3723 5918 4021 5924
rect 3708 5326 3747 5807
rect 3190 5287 3747 5326
rect 3819 5328 3858 5738
rect 4217 5653 4261 6422
rect 4331 6265 4362 6475
rect 4421 6157 4521 6415
rect 4339 6151 4637 6157
rect 4339 5924 4351 6151
rect 4625 5924 4637 6151
rect 4339 5918 4637 5924
rect 4324 5328 4363 5807
rect 3819 5289 4363 5328
rect 4445 5328 4484 5745
rect 4833 5653 4877 6422
rect 4947 6265 4978 6475
rect 5037 6157 5137 6415
rect 4955 6151 5253 6157
rect 4955 5924 4967 6151
rect 5241 5924 5253 6151
rect 4955 5918 5253 5924
rect 4940 5328 4979 5807
rect 4445 5289 4979 5328
rect 5048 5328 5087 5737
rect 5449 5653 5493 6422
rect 5563 6265 5594 6475
rect 5653 6157 5753 6415
rect 5872 6338 5923 6475
rect 6078 6159 6178 6421
rect 6386 6173 6396 6272
rect 6756 6173 6766 6272
rect 5571 6151 5869 6157
rect 5571 5924 5583 6151
rect 5857 5924 5869 6151
rect 5571 5918 5869 5924
rect 6069 6150 6246 6159
rect 6069 5924 6077 6150
rect 6236 5924 6246 6150
rect 6069 5917 6246 5924
rect 5556 5328 5595 5807
rect 5672 5332 5711 5744
rect 6395 5666 6479 6173
rect 6904 5967 6914 5988
rect 5048 5289 5595 5328
rect 3060 5163 3070 5286
rect 2472 5026 2482 5088
rect 2639 5026 2649 5088
rect 2459 4752 2496 4959
rect 2180 4715 2496 4752
rect 2205 4605 2484 4611
rect 2205 4448 2217 4605
rect 2472 4448 2484 4605
rect 2205 4442 2484 4448
rect 2303 4431 2395 4442
rect 2311 4188 2395 4431
rect 2461 4130 2494 4333
rect 2561 4188 2603 4877
rect 2904 4681 2946 4874
rect 3016 4720 3055 5163
rect 3190 5015 3229 5287
rect 3128 4976 3229 5015
rect 3128 4787 3167 4976
rect 3460 4681 3502 4874
rect 3572 4720 3611 5287
rect 3819 5016 3858 5289
rect 3679 4977 3858 5016
rect 3679 4781 3718 4977
rect 4016 4681 4058 4874
rect 4128 4720 4167 5289
rect 4445 5018 4484 5289
rect 4235 4979 4484 5018
rect 4235 4789 4274 4979
rect 4572 4681 4614 4874
rect 4684 4720 4723 5289
rect 5048 5021 5087 5289
rect 4789 4982 5087 5021
rect 4789 4781 4828 4982
rect 5128 4681 5170 4874
rect 5240 4720 5279 5289
rect 5659 5167 5669 5332
rect 5726 5290 5736 5332
rect 6540 5290 6584 5941
rect 5726 5223 6584 5290
rect 6642 5929 6914 5967
rect 5726 5167 5736 5223
rect 5672 5020 5711 5167
rect 5347 4981 5711 5020
rect 5347 4782 5386 4981
rect 2904 4639 3159 4681
rect 3460 4639 3715 4681
rect 4016 4639 4271 4681
rect 4572 4639 4827 4681
rect 5128 4639 5383 4681
rect 2761 4605 3040 4611
rect 2761 4448 2773 4605
rect 3028 4448 3040 4605
rect 2761 4442 3040 4448
rect 2859 4431 2951 4442
rect 2867 4188 2951 4431
rect 3017 4130 3050 4333
rect 3117 4188 3159 4639
rect 3317 4605 3596 4611
rect 3317 4448 3329 4605
rect 3584 4448 3596 4605
rect 3317 4442 3596 4448
rect 3415 4431 3507 4442
rect 3423 4188 3507 4431
rect 3573 4130 3606 4333
rect 3673 4188 3715 4639
rect 3873 4605 4152 4611
rect 3873 4448 3885 4605
rect 4140 4448 4152 4605
rect 3873 4442 4152 4448
rect 3971 4431 4063 4442
rect 3979 4188 4063 4431
rect 4129 4130 4162 4333
rect 4229 4188 4271 4639
rect 4429 4605 4708 4611
rect 4429 4448 4441 4605
rect 4696 4448 4708 4605
rect 4429 4442 4708 4448
rect 4527 4431 4619 4442
rect 4535 4188 4619 4431
rect 4685 4130 4718 4333
rect 4785 4188 4827 4639
rect 4985 4605 5264 4611
rect 4985 4448 4997 4605
rect 5252 4448 5264 4605
rect 4985 4442 5264 4448
rect 5083 4431 5175 4442
rect 5091 4188 5175 4431
rect 5241 4130 5274 4333
rect 5341 4188 5383 4639
rect 5674 4618 5842 4630
rect 5674 4613 5680 4618
rect 5540 4605 5680 4613
rect 5540 4448 5549 4605
rect 5836 4449 5842 4618
rect 5804 4448 5842 4449
rect 5540 4439 5842 4448
rect 5674 4437 5842 4439
rect 6087 4447 6131 5223
rect 6428 4623 6466 4860
rect 6533 4743 6569 4933
rect 6642 4785 6680 5929
rect 6904 5910 6914 5929
rect 7105 5910 7115 5988
rect 6934 5145 7307 5179
rect 6934 4961 6968 5145
rect 6814 4897 6824 4961
rect 7011 4897 7021 4961
rect 6533 4707 6956 4743
rect 6917 4638 6956 4707
rect 6428 4585 6679 4623
rect 6917 4599 6981 4638
rect 5708 4274 5792 4437
rect 6087 4404 6574 4447
rect 6218 4403 6574 4404
rect 5708 4273 6468 4274
rect 5708 4191 6478 4273
rect 5708 4190 6366 4191
rect 1454 4081 5518 4129
rect 6530 4124 6574 4403
rect 6641 4190 6679 4585
rect 6971 4574 6981 4599
rect 7168 4574 7178 4638
rect 8721 4316 8764 6841
rect 8609 4306 8764 4316
rect 7152 4256 8764 4306
rect 106 3993 199 4005
rect 1129 3928 6787 4013
rect 1129 3873 1183 3928
rect 6742 3873 6787 3928
rect 7152 3923 7196 4256
rect 8600 3943 8764 4256
rect 8829 6801 8915 6841
rect 10141 6801 10178 6866
rect 8829 6774 10178 6801
rect 8829 3943 8898 6774
rect 10302 6702 10377 7607
rect 9378 6627 10377 6702
rect 9151 6483 9161 6555
rect 9337 6483 9347 6555
rect 9138 5988 9191 6188
rect 9275 6102 9337 6483
rect 8949 5916 8959 5988
rect 9135 5934 9191 5988
rect 9135 5916 9145 5934
rect 9236 5780 9268 6064
rect 9124 5708 9134 5780
rect 9310 5708 9320 5780
rect 9236 5641 9268 5643
rect 9096 5569 9106 5641
rect 9282 5569 9292 5641
rect 9378 4131 9453 6627
rect 9505 6573 9825 6579
rect 9505 6444 9517 6573
rect 9813 6444 9825 6573
rect 10508 6564 10886 7121
rect 9505 6438 9825 6444
rect 10026 6554 10886 6564
rect 10026 6455 10037 6554
rect 10397 6455 10886 6554
rect 10026 6364 10886 6455
rect 9522 6177 9532 6276
rect 9892 6177 9902 6276
rect 10026 6249 10723 6364
rect 9528 4934 9690 6177
rect 10026 6122 10507 6249
rect 10711 6122 10723 6249
rect 10026 6116 10723 6122
rect 10026 6039 10615 6116
rect 10026 6023 10722 6039
rect 10026 5960 10500 6023
rect 10607 5960 10722 6023
rect 10822 5989 10870 6044
rect 10026 5945 10722 5960
rect 10026 5943 10226 5945
rect 10713 5944 10722 5945
rect 10702 5829 10788 5883
rect 10702 5672 10743 5829
rect 10820 5782 10870 5989
rect 10373 5655 10383 5672
rect 10312 5600 10383 5655
rect 10559 5614 10743 5672
rect 10559 5600 10569 5614
rect 10312 5290 10350 5600
rect 10633 5581 10699 5614
rect 10771 5613 10781 5782
rect 10850 5622 10870 5782
rect 10850 5613 10860 5622
rect 10479 5388 10599 5400
rect 10222 5252 10350 5290
rect 10222 5136 10260 5252
rect 10387 5222 10485 5388
rect 10319 5192 10485 5222
rect 10521 5192 10599 5388
rect 10819 5211 10860 5613
rect 10319 5140 10599 5192
rect 10137 5026 10147 5098
rect 10323 5026 10333 5098
rect 10387 4934 10599 5140
rect 10744 4950 10780 5135
rect 9528 4734 10599 4934
rect 10661 4891 10671 4950
rect 10857 4891 10867 4950
rect 10039 4680 10599 4734
rect 10039 4191 10886 4680
rect 9378 4056 10397 4131
rect 8600 3923 8898 3943
rect 7152 3892 8898 3923
rect 1129 3856 6787 3873
rect 1850 3768 3533 3774
rect 1850 3689 1862 3768
rect 3521 3689 3533 3768
rect 1850 3683 3533 3689
rect 5362 3771 7045 3777
rect 5362 3692 5374 3771
rect 7033 3692 7045 3771
rect 5362 3686 7045 3692
rect 86 3543 605 3550
rect 86 3134 100 3543
rect 351 3134 605 3543
rect 86 3118 605 3134
rect 700 3118 936 3550
rect 1032 3118 1268 3550
rect 1364 3118 1600 3550
rect 1696 3118 1932 3550
rect 2028 3118 2264 3550
rect 2360 3118 2596 3550
rect 2692 3118 2928 3550
rect 3024 3118 3260 3550
rect 3356 3118 3592 3550
rect 3688 3118 3924 3550
rect 4020 3118 4256 3550
rect 4352 3118 4588 3550
rect 4684 3118 4920 3550
rect 5016 3118 5252 3550
rect 5348 3118 5584 3550
rect 5680 3118 5916 3550
rect 6012 3118 6248 3550
rect 6344 3118 6580 3550
rect 6676 3118 6912 3550
rect 7008 3118 7244 3550
rect 7340 3118 7576 3550
rect 7672 3118 7908 3550
rect 8004 3118 8240 3550
rect 8336 3118 8572 3550
rect 8668 3118 8904 3550
rect 9000 3118 9236 3550
rect 9332 3118 9568 3550
rect 9664 3118 9900 3550
rect 9996 3118 10232 3550
rect 10322 3115 10397 4056
rect 10508 3634 10886 4191
rect 313 3045 419 3057
rect 10478 3046 10584 3058
rect 309 1960 319 3045
rect 413 1960 423 3045
rect 10474 1961 10484 3046
rect 10578 1961 10588 3046
rect 313 1948 419 1960
rect 10478 1949 10584 1961
rect 534 1218 770 1650
rect 866 1218 1102 1650
rect 1198 1218 1434 1650
rect 1530 1218 1766 1650
rect 1862 1218 2098 1650
rect 2194 1218 2430 1650
rect 2526 1218 2762 1650
rect 2858 1218 3094 1650
rect 3190 1218 3426 1650
rect 3522 1218 3758 1650
rect 3854 1218 4090 1650
rect 4186 1218 4422 1650
rect 4518 1218 4754 1650
rect 4850 1218 5086 1650
rect 5182 1218 5418 1650
rect 5514 1218 5750 1650
rect 5846 1218 6082 1650
rect 6178 1218 6414 1650
rect 6510 1218 6746 1650
rect 6842 1218 7078 1650
rect 7174 1218 7410 1650
rect 7506 1218 7742 1650
rect 7838 1218 8074 1650
rect 8170 1218 8406 1650
rect 8502 1218 8738 1650
rect 8834 1218 9070 1650
rect 9166 1218 9402 1650
rect 9498 1218 9734 1650
rect 9830 1218 10066 1650
rect 10162 1218 10398 1650
<< via1 >>
rect 10698 7712 10786 8810
rect 112 4005 193 7683
rect 654 6942 1795 7069
rect 8761 6901 10142 6999
rect 2190 6753 6770 6818
rect 7203 6547 8607 6880
rect 2503 5924 2777 6151
rect 1449 4905 1606 4967
rect 1122 4442 1278 4611
rect 1970 5022 2127 5084
rect 1661 4448 1916 4605
rect 3119 5924 3393 6151
rect 3003 5163 3060 5328
rect 3735 5924 4009 6151
rect 4351 5924 4625 6151
rect 4967 5924 5241 6151
rect 6396 6173 6756 6272
rect 5583 5924 5857 6151
rect 6077 5924 6236 6150
rect 2482 5026 2639 5088
rect 2217 4448 2472 4605
rect 5669 5167 5726 5332
rect 2773 4448 3028 4605
rect 3329 4448 3584 4605
rect 3885 4448 4140 4605
rect 4441 4448 4696 4605
rect 4997 4448 5252 4605
rect 5549 4449 5680 4605
rect 5680 4449 5804 4605
rect 5549 4448 5804 4449
rect 6914 5910 7105 5988
rect 6824 4897 7011 4961
rect 6981 4574 7168 4638
rect 1183 3873 6742 3928
rect 7196 3923 8600 4256
rect 9161 6483 9337 6555
rect 8959 5916 9135 5988
rect 9134 5708 9310 5780
rect 9106 5569 9282 5641
rect 9517 6444 9813 6573
rect 10037 6455 10397 6554
rect 9532 6177 9892 6276
rect 10383 5600 10559 5672
rect 10781 5613 10850 5782
rect 9871 5022 9930 5208
rect 10147 5026 10323 5098
rect 10671 4891 10857 4950
rect 1862 3689 3521 3768
rect 5374 3692 7033 3771
rect 100 3134 351 3543
rect 319 1960 413 3045
rect 10484 1961 10578 3046
<< metal2 >>
rect 10698 8819 10786 8820
rect 0 8810 10886 8819
rect 0 7712 10698 8810
rect 10786 7712 10886 8810
rect 0 7701 10886 7712
rect 92 7683 358 7701
rect 92 4005 112 7683
rect 193 4005 358 7683
rect 627 7069 1828 7083
rect 627 7065 654 7069
rect 92 3543 358 4005
rect 92 3134 100 3543
rect 351 3134 358 3543
rect 92 3128 358 3134
rect 625 6942 654 7065
rect 1795 6942 1828 7069
rect 625 6925 1828 6942
rect 625 6878 1175 6925
rect 625 5294 1174 6878
rect 2453 6865 4111 7701
rect 5409 6865 7067 7701
rect 9837 7156 10178 7701
rect 7169 6901 8652 7090
rect 8721 6999 10178 7156
rect 8721 6901 8761 6999
rect 10142 6901 10178 6999
rect 7169 6880 8651 6901
rect 8721 6882 10178 6901
rect 2119 6818 6838 6865
rect 2119 6753 2190 6818
rect 6770 6753 6838 6818
rect 2119 6655 6838 6753
rect 2453 6199 4111 6655
rect 5409 6199 5951 6655
rect 7169 6547 7203 6880
rect 8607 6547 8651 6880
rect 9517 6574 9813 6583
rect 7169 6506 8651 6547
rect 9147 6573 10402 6574
rect 9147 6555 9517 6573
rect 9147 6483 9161 6555
rect 9337 6483 9517 6555
rect 9147 6444 9517 6483
rect 9813 6554 10402 6573
rect 9813 6455 10037 6554
rect 10397 6455 10402 6554
rect 9813 6444 10402 6455
rect 9147 6442 10402 6444
rect 9517 6434 9813 6442
rect 6396 6274 6756 6282
rect 9532 6276 9892 6286
rect 6396 6272 9532 6274
rect 1538 6151 6284 6199
rect 6756 6177 9532 6272
rect 6756 6176 9892 6177
rect 6396 6163 6756 6173
rect 9532 6167 9892 6176
rect 1538 5924 2503 6151
rect 2777 5924 3119 6151
rect 3393 5924 3735 6151
rect 4009 5924 4351 6151
rect 4625 5924 4967 6151
rect 5241 5924 5583 6151
rect 5857 6150 6284 6151
rect 5857 5924 6077 6150
rect 6236 5924 6284 6150
rect 1538 5883 6284 5924
rect 6914 5988 7105 5998
rect 8959 5988 9135 5998
rect 7105 5929 8856 5973
rect 8958 5929 8959 5973
rect 6914 5900 7105 5910
rect 8812 5876 8856 5929
rect 10770 5973 10970 6050
rect 9135 5929 10970 5973
rect 8959 5906 9135 5916
rect 8812 5832 10308 5876
rect 10770 5850 10970 5929
rect 9134 5780 9310 5790
rect 9134 5698 9310 5708
rect 10264 5654 10308 5832
rect 10781 5782 10850 5850
rect 10383 5672 10559 5682
rect 9106 5641 9282 5651
rect 3003 5328 3060 5338
rect 625 4644 1175 5294
rect 5669 5332 5726 5342
rect 3060 5220 5669 5261
rect 3003 5153 3060 5163
rect 5669 5157 5726 5167
rect 1970 5084 2127 5094
rect 2482 5088 2639 5098
rect 1932 5023 1970 5084
rect 2127 5026 2482 5084
rect 2639 5026 7147 5084
rect 2127 5023 7147 5026
rect 1970 5012 2127 5022
rect 2482 5016 2639 5023
rect 1449 4967 1606 4977
rect 6814 4961 7011 4971
rect 6814 4950 6824 4961
rect 1606 4905 6824 4950
rect 1449 4895 1606 4905
rect 6824 4887 7011 4897
rect 7086 4926 7147 5023
rect 7086 4865 7916 4926
rect 625 4611 6019 4644
rect 6981 4639 7168 4648
rect 8572 4639 8637 5600
rect 10264 5610 10383 5654
rect 10781 5603 10850 5613
rect 10383 5590 10559 5600
rect 9106 5559 9282 5569
rect 9900 5391 10453 5445
rect 9863 5022 9871 5208
rect 9930 5022 9939 5208
rect 10147 5098 10323 5108
rect 10399 5086 10453 5391
rect 10323 5053 10453 5086
rect 10770 5053 10970 5196
rect 10323 5039 10970 5053
rect 9871 4951 9930 5022
rect 10147 5016 10323 5026
rect 10399 4999 10970 5039
rect 10770 4996 10970 4999
rect 10671 4951 10857 4958
rect 9871 4950 10857 4951
rect 9871 4892 10671 4950
rect 10671 4881 10857 4891
rect 625 4442 1122 4611
rect 1278 4605 6019 4611
rect 1278 4448 1661 4605
rect 1916 4448 2217 4605
rect 2472 4448 2773 4605
rect 3028 4448 3329 4605
rect 3584 4448 3885 4605
rect 4140 4448 4441 4605
rect 4696 4448 4997 4605
rect 5252 4448 5549 4605
rect 5804 4448 6019 4605
rect 6979 4638 8637 4639
rect 6979 4574 6981 4638
rect 7168 4574 8637 4638
rect 6981 4564 7168 4574
rect 1278 4442 6019 4448
rect 625 4342 6019 4442
rect 625 4038 1175 4342
rect 1861 4038 3520 4342
rect 5375 4038 5918 4342
rect 7152 4256 8634 4306
rect 625 3928 6814 4038
rect 625 3873 1183 3928
rect 6742 3873 6814 3928
rect 7152 3923 7196 4256
rect 8600 3923 8634 4256
rect 7152 3892 8634 3923
rect 625 3824 6814 3873
rect 625 3062 1175 3824
rect 1861 3768 3521 3824
rect 1861 3689 1862 3768
rect 1861 3679 3521 3689
rect 5374 3771 7034 3824
rect 7033 3692 7034 3771
rect 5374 3682 7034 3692
rect 1861 3062 3520 3679
rect 5375 3062 7034 3682
rect 0 3046 10886 3062
rect 0 3045 10484 3046
rect 0 1960 319 3045
rect 413 1961 10484 3045
rect 10578 1961 10886 3046
rect 413 1960 10886 1961
rect 0 1944 10886 1960
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D3 paramcells
timestamp 1699295625
transform 1 0 9223 0 1 5604
box -183 -183 183 183
use level_shifter  level_shifter_0
timestamp 1699295625
transform -1 0 9816 0 -1 4214
box -422 -2544 2736 144
use sky130_fd_pr__nfet_01v8_L9WNCD  sky130_fd_pr__nfet_01v8_L9WNCD_0 paramcells
timestamp 1699295625
transform 1 0 10759 0 1 5958
box -211 -229 211 229
use sky130_fd_pr__pfet_01v8_2Z69BZ  sky130_fd_pr__pfet_01v8_2Z69BZ_0 paramcells
timestamp 1699295625
transform 1 0 10286 0 1 5145
box -211 -226 211 226
use sky130_fd_pr__pfet_01v8_856REK  sky130_fd_pr__pfet_01v8_856REK_0 paramcells
timestamp 1716055179
transform 1 0 10714 0 -1 5350
box -263 -369 263 369
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  sky130_fd_pr__pfet_g5v0d10v5_6ELFTH_0 paramcells
timestamp 1699295625
transform 1 0 2498 0 1 6373
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  sky130_fd_pr__pfet_g5v0d10v5_6ELFTH_1
timestamp 1699295625
transform 1 0 1646 0 1 6373
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  sky130_fd_pr__pfet_g5v0d10v5_6ELFTH_2
timestamp 1699295625
transform 1 0 2072 0 1 6373
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  sky130_fd_pr__pfet_g5v0d10v5_6ELFTH_3
timestamp 1699295625
transform 1 0 2498 0 1 5695
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  sky130_fd_pr__pfet_g5v0d10v5_6ELFTH_4
timestamp 1699295625
transform 1 0 2072 0 1 5695
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  sky130_fd_pr__pfet_g5v0d10v5_6ELFTH_5
timestamp 1699295625
transform 1 0 5578 0 1 6373
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_T537S5  sky130_fd_pr__pfet_g5v0d10v5_T537S5_0 paramcells
timestamp 1716055179
transform 1 0 6560 0 1 5752
box -308 -423 308 423
use sky130_fd_pr__res_xhigh_po_0p35_NVJ5PF  sky130_fd_pr__res_xhigh_po_0p35_NVJ5PF_0 paramcells
timestamp 1715996061
transform 1 0 5466 0 1 2384
box -5098 -1332 5098 1332
use sky130_fd_pr__res_xhigh_po_0p35_NVJ5PF  sky130_fd_pr__res_xhigh_po_0p35_NVJ5PF_1
timestamp 1715996061
transform 1 0 5446 0 1 8334
box -5098 -1332 5098 1332
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM1 paramcells
timestamp 1699295625
transform 1 0 3032 0 1 4830
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM2
timestamp 1699295625
transform 1 0 3114 0 1 5695
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM3
timestamp 1699295625
transform 1 0 3730 0 1 5695
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM4
timestamp 1699295625
transform 1 0 3588 0 1 4830
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM7
timestamp 1699295625
transform 1 0 4962 0 1 5695
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM8
timestamp 1699295625
transform 1 0 4700 0 1 4830
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM9
timestamp 1699295625
transform 1 0 4346 0 1 5695
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM10
timestamp 1699295625
transform 1 0 4144 0 1 4830
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM12
timestamp 1699295625
transform 1 0 6552 0 1 4228
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM13
timestamp 1699295625
transform 1 0 6552 0 1 4828
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM15
timestamp 1699295625
transform 1 0 5578 0 1 5695
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM16
timestamp 1699295625
transform 1 0 5256 0 1 4830
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM17
timestamp 1699295625
transform 1 0 4962 0 1 6373
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM18
timestamp 1699295625
transform 1 0 6004 0 1 6373
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM19
timestamp 1699295625
transform 1 0 5256 0 1 4230
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM20
timestamp 1699295625
transform 1 0 4700 0 1 4230
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM21
timestamp 1699295625
transform 1 0 1920 0 1 4230
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM23
timestamp 1699295625
transform 1 0 1920 0 1 4828
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM24
timestamp 1699295625
transform 1 0 3114 0 1 6373
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM25
timestamp 1699295625
transform 1 0 3730 0 1 6373
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM26
timestamp 1699295625
transform 1 0 4346 0 1 6373
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM27
timestamp 1699295625
transform 1 0 4144 0 1 4230
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM28
timestamp 1699295625
transform 1 0 3588 0 1 4230
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM29
timestamp 1699295625
transform 1 0 3032 0 1 4230
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM30
timestamp 1699295625
transform 1 0 2476 0 1 4230
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM33
timestamp 1699295625
transform 1 0 1364 0 1 4828
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM34
timestamp 1699295625
transform 1 0 1646 0 1 5695
box -308 -339 308 339
use sky130_fd_pr__nfet_01v8_L7BSKG  XM35 paramcells
timestamp 1699295625
transform 1 0 9251 0 1 6113
box -211 -221 211 221
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM36
timestamp 1699295625
transform 1 0 2476 0 1 4830
box -278 -300 278 300
<< labels >>
flabel metal2 0 7701 200 8819 0 FreeSans 256 0 0 0 avdd
port 0 nsew
flabel metal2 0 1944 200 3062 0 FreeSans 256 0 0 0 avss
port 1 nsew
flabel metal2 s 10786 7701 10886 8819 0 FreeSans 640 90 0 0 avdd
port 0 nsew
flabel metal1 10686 6364 10886 7121 0 FreeSans 256 0 0 0 dvss
port 2 nsew
flabel metal2 s 10578 1944 10886 3062 0 FreeSans 960 90 0 0 avss
port 1 nsew
flabel metal1 10686 3634 10886 4391 0 FreeSans 256 0 0 0 dvdd
port 3 nsew
flabel metal2 10770 5850 10970 6050 0 FreeSans 256 0 0 0 dout
port 5 nsew
flabel metal2 10770 4996 10970 5196 0 FreeSans 256 0 0 0 ena
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 12242 10724
<< end >>
