magic
tech sky130A
magscale 1 2
timestamp 1715996061
<< pwell >>
rect -5098 -1332 5098 1332
<< psubdiff >>
rect -5062 1262 -4966 1296
rect 4966 1262 5062 1296
rect -5062 1200 -5028 1262
rect 5028 1200 5062 1262
rect -5062 -1262 -5028 -1200
rect 5028 -1262 5062 -1200
rect -5062 -1296 -4966 -1262
rect 4966 -1296 5062 -1262
<< psubdiffcont >>
rect -4966 1262 4966 1296
rect -5062 -1200 -5028 1200
rect 5028 -1200 5062 1200
rect -4966 -1296 4966 -1262
<< xpolycontact >>
rect -4932 734 -4862 1166
rect -4932 -1166 -4862 -734
rect -4766 734 -4696 1166
rect -4766 -1166 -4696 -734
rect -4600 734 -4530 1166
rect -4600 -1166 -4530 -734
rect -4434 734 -4364 1166
rect -4434 -1166 -4364 -734
rect -4268 734 -4198 1166
rect -4268 -1166 -4198 -734
rect -4102 734 -4032 1166
rect -4102 -1166 -4032 -734
rect -3936 734 -3866 1166
rect -3936 -1166 -3866 -734
rect -3770 734 -3700 1166
rect -3770 -1166 -3700 -734
rect -3604 734 -3534 1166
rect -3604 -1166 -3534 -734
rect -3438 734 -3368 1166
rect -3438 -1166 -3368 -734
rect -3272 734 -3202 1166
rect -3272 -1166 -3202 -734
rect -3106 734 -3036 1166
rect -3106 -1166 -3036 -734
rect -2940 734 -2870 1166
rect -2940 -1166 -2870 -734
rect -2774 734 -2704 1166
rect -2774 -1166 -2704 -734
rect -2608 734 -2538 1166
rect -2608 -1166 -2538 -734
rect -2442 734 -2372 1166
rect -2442 -1166 -2372 -734
rect -2276 734 -2206 1166
rect -2276 -1166 -2206 -734
rect -2110 734 -2040 1166
rect -2110 -1166 -2040 -734
rect -1944 734 -1874 1166
rect -1944 -1166 -1874 -734
rect -1778 734 -1708 1166
rect -1778 -1166 -1708 -734
rect -1612 734 -1542 1166
rect -1612 -1166 -1542 -734
rect -1446 734 -1376 1166
rect -1446 -1166 -1376 -734
rect -1280 734 -1210 1166
rect -1280 -1166 -1210 -734
rect -1114 734 -1044 1166
rect -1114 -1166 -1044 -734
rect -948 734 -878 1166
rect -948 -1166 -878 -734
rect -782 734 -712 1166
rect -782 -1166 -712 -734
rect -616 734 -546 1166
rect -616 -1166 -546 -734
rect -450 734 -380 1166
rect -450 -1166 -380 -734
rect -284 734 -214 1166
rect -284 -1166 -214 -734
rect -118 734 -48 1166
rect -118 -1166 -48 -734
rect 48 734 118 1166
rect 48 -1166 118 -734
rect 214 734 284 1166
rect 214 -1166 284 -734
rect 380 734 450 1166
rect 380 -1166 450 -734
rect 546 734 616 1166
rect 546 -1166 616 -734
rect 712 734 782 1166
rect 712 -1166 782 -734
rect 878 734 948 1166
rect 878 -1166 948 -734
rect 1044 734 1114 1166
rect 1044 -1166 1114 -734
rect 1210 734 1280 1166
rect 1210 -1166 1280 -734
rect 1376 734 1446 1166
rect 1376 -1166 1446 -734
rect 1542 734 1612 1166
rect 1542 -1166 1612 -734
rect 1708 734 1778 1166
rect 1708 -1166 1778 -734
rect 1874 734 1944 1166
rect 1874 -1166 1944 -734
rect 2040 734 2110 1166
rect 2040 -1166 2110 -734
rect 2206 734 2276 1166
rect 2206 -1166 2276 -734
rect 2372 734 2442 1166
rect 2372 -1166 2442 -734
rect 2538 734 2608 1166
rect 2538 -1166 2608 -734
rect 2704 734 2774 1166
rect 2704 -1166 2774 -734
rect 2870 734 2940 1166
rect 2870 -1166 2940 -734
rect 3036 734 3106 1166
rect 3036 -1166 3106 -734
rect 3202 734 3272 1166
rect 3202 -1166 3272 -734
rect 3368 734 3438 1166
rect 3368 -1166 3438 -734
rect 3534 734 3604 1166
rect 3534 -1166 3604 -734
rect 3700 734 3770 1166
rect 3700 -1166 3770 -734
rect 3866 734 3936 1166
rect 3866 -1166 3936 -734
rect 4032 734 4102 1166
rect 4032 -1166 4102 -734
rect 4198 734 4268 1166
rect 4198 -1166 4268 -734
rect 4364 734 4434 1166
rect 4364 -1166 4434 -734
rect 4530 734 4600 1166
rect 4530 -1166 4600 -734
rect 4696 734 4766 1166
rect 4696 -1166 4766 -734
rect 4862 734 4932 1166
rect 4862 -1166 4932 -734
<< xpolyres >>
rect -4932 -734 -4862 734
rect -4766 -734 -4696 734
rect -4600 -734 -4530 734
rect -4434 -734 -4364 734
rect -4268 -734 -4198 734
rect -4102 -734 -4032 734
rect -3936 -734 -3866 734
rect -3770 -734 -3700 734
rect -3604 -734 -3534 734
rect -3438 -734 -3368 734
rect -3272 -734 -3202 734
rect -3106 -734 -3036 734
rect -2940 -734 -2870 734
rect -2774 -734 -2704 734
rect -2608 -734 -2538 734
rect -2442 -734 -2372 734
rect -2276 -734 -2206 734
rect -2110 -734 -2040 734
rect -1944 -734 -1874 734
rect -1778 -734 -1708 734
rect -1612 -734 -1542 734
rect -1446 -734 -1376 734
rect -1280 -734 -1210 734
rect -1114 -734 -1044 734
rect -948 -734 -878 734
rect -782 -734 -712 734
rect -616 -734 -546 734
rect -450 -734 -380 734
rect -284 -734 -214 734
rect -118 -734 -48 734
rect 48 -734 118 734
rect 214 -734 284 734
rect 380 -734 450 734
rect 546 -734 616 734
rect 712 -734 782 734
rect 878 -734 948 734
rect 1044 -734 1114 734
rect 1210 -734 1280 734
rect 1376 -734 1446 734
rect 1542 -734 1612 734
rect 1708 -734 1778 734
rect 1874 -734 1944 734
rect 2040 -734 2110 734
rect 2206 -734 2276 734
rect 2372 -734 2442 734
rect 2538 -734 2608 734
rect 2704 -734 2774 734
rect 2870 -734 2940 734
rect 3036 -734 3106 734
rect 3202 -734 3272 734
rect 3368 -734 3438 734
rect 3534 -734 3604 734
rect 3700 -734 3770 734
rect 3866 -734 3936 734
rect 4032 -734 4102 734
rect 4198 -734 4268 734
rect 4364 -734 4434 734
rect 4530 -734 4600 734
rect 4696 -734 4766 734
rect 4862 -734 4932 734
<< locali >>
rect -5062 1262 -4966 1296
rect 4966 1262 5062 1296
rect -5062 1200 -5028 1262
rect 5028 1200 5062 1262
rect -5062 -1262 -5028 -1200
rect 5028 -1262 5062 -1200
rect -5062 -1296 -4966 -1262
rect 4966 -1296 5062 -1262
<< viali >>
rect -4916 751 -4878 1148
rect -4750 751 -4712 1148
rect -4584 751 -4546 1148
rect -4418 751 -4380 1148
rect -4252 751 -4214 1148
rect -4086 751 -4048 1148
rect -3920 751 -3882 1148
rect -3754 751 -3716 1148
rect -3588 751 -3550 1148
rect -3422 751 -3384 1148
rect -3256 751 -3218 1148
rect -3090 751 -3052 1148
rect -2924 751 -2886 1148
rect -2758 751 -2720 1148
rect -2592 751 -2554 1148
rect -2426 751 -2388 1148
rect -2260 751 -2222 1148
rect -2094 751 -2056 1148
rect -1928 751 -1890 1148
rect -1762 751 -1724 1148
rect -1596 751 -1558 1148
rect -1430 751 -1392 1148
rect -1264 751 -1226 1148
rect -1098 751 -1060 1148
rect -932 751 -894 1148
rect -766 751 -728 1148
rect -600 751 -562 1148
rect -434 751 -396 1148
rect -268 751 -230 1148
rect -102 751 -64 1148
rect 64 751 102 1148
rect 230 751 268 1148
rect 396 751 434 1148
rect 562 751 600 1148
rect 728 751 766 1148
rect 894 751 932 1148
rect 1060 751 1098 1148
rect 1226 751 1264 1148
rect 1392 751 1430 1148
rect 1558 751 1596 1148
rect 1724 751 1762 1148
rect 1890 751 1928 1148
rect 2056 751 2094 1148
rect 2222 751 2260 1148
rect 2388 751 2426 1148
rect 2554 751 2592 1148
rect 2720 751 2758 1148
rect 2886 751 2924 1148
rect 3052 751 3090 1148
rect 3218 751 3256 1148
rect 3384 751 3422 1148
rect 3550 751 3588 1148
rect 3716 751 3754 1148
rect 3882 751 3920 1148
rect 4048 751 4086 1148
rect 4214 751 4252 1148
rect 4380 751 4418 1148
rect 4546 751 4584 1148
rect 4712 751 4750 1148
rect 4878 751 4916 1148
rect -4916 -1148 -4878 -751
rect -4750 -1148 -4712 -751
rect -4584 -1148 -4546 -751
rect -4418 -1148 -4380 -751
rect -4252 -1148 -4214 -751
rect -4086 -1148 -4048 -751
rect -3920 -1148 -3882 -751
rect -3754 -1148 -3716 -751
rect -3588 -1148 -3550 -751
rect -3422 -1148 -3384 -751
rect -3256 -1148 -3218 -751
rect -3090 -1148 -3052 -751
rect -2924 -1148 -2886 -751
rect -2758 -1148 -2720 -751
rect -2592 -1148 -2554 -751
rect -2426 -1148 -2388 -751
rect -2260 -1148 -2222 -751
rect -2094 -1148 -2056 -751
rect -1928 -1148 -1890 -751
rect -1762 -1148 -1724 -751
rect -1596 -1148 -1558 -751
rect -1430 -1148 -1392 -751
rect -1264 -1148 -1226 -751
rect -1098 -1148 -1060 -751
rect -932 -1148 -894 -751
rect -766 -1148 -728 -751
rect -600 -1148 -562 -751
rect -434 -1148 -396 -751
rect -268 -1148 -230 -751
rect -102 -1148 -64 -751
rect 64 -1148 102 -751
rect 230 -1148 268 -751
rect 396 -1148 434 -751
rect 562 -1148 600 -751
rect 728 -1148 766 -751
rect 894 -1148 932 -751
rect 1060 -1148 1098 -751
rect 1226 -1148 1264 -751
rect 1392 -1148 1430 -751
rect 1558 -1148 1596 -751
rect 1724 -1148 1762 -751
rect 1890 -1148 1928 -751
rect 2056 -1148 2094 -751
rect 2222 -1148 2260 -751
rect 2388 -1148 2426 -751
rect 2554 -1148 2592 -751
rect 2720 -1148 2758 -751
rect 2886 -1148 2924 -751
rect 3052 -1148 3090 -751
rect 3218 -1148 3256 -751
rect 3384 -1148 3422 -751
rect 3550 -1148 3588 -751
rect 3716 -1148 3754 -751
rect 3882 -1148 3920 -751
rect 4048 -1148 4086 -751
rect 4214 -1148 4252 -751
rect 4380 -1148 4418 -751
rect 4546 -1148 4584 -751
rect 4712 -1148 4750 -751
rect 4878 -1148 4916 -751
<< metal1 >>
rect -4922 1148 -4872 1160
rect -4922 751 -4916 1148
rect -4878 751 -4872 1148
rect -4922 739 -4872 751
rect -4756 1148 -4706 1160
rect -4756 751 -4750 1148
rect -4712 751 -4706 1148
rect -4756 739 -4706 751
rect -4590 1148 -4540 1160
rect -4590 751 -4584 1148
rect -4546 751 -4540 1148
rect -4590 739 -4540 751
rect -4424 1148 -4374 1160
rect -4424 751 -4418 1148
rect -4380 751 -4374 1148
rect -4424 739 -4374 751
rect -4258 1148 -4208 1160
rect -4258 751 -4252 1148
rect -4214 751 -4208 1148
rect -4258 739 -4208 751
rect -4092 1148 -4042 1160
rect -4092 751 -4086 1148
rect -4048 751 -4042 1148
rect -4092 739 -4042 751
rect -3926 1148 -3876 1160
rect -3926 751 -3920 1148
rect -3882 751 -3876 1148
rect -3926 739 -3876 751
rect -3760 1148 -3710 1160
rect -3760 751 -3754 1148
rect -3716 751 -3710 1148
rect -3760 739 -3710 751
rect -3594 1148 -3544 1160
rect -3594 751 -3588 1148
rect -3550 751 -3544 1148
rect -3594 739 -3544 751
rect -3428 1148 -3378 1160
rect -3428 751 -3422 1148
rect -3384 751 -3378 1148
rect -3428 739 -3378 751
rect -3262 1148 -3212 1160
rect -3262 751 -3256 1148
rect -3218 751 -3212 1148
rect -3262 739 -3212 751
rect -3096 1148 -3046 1160
rect -3096 751 -3090 1148
rect -3052 751 -3046 1148
rect -3096 739 -3046 751
rect -2930 1148 -2880 1160
rect -2930 751 -2924 1148
rect -2886 751 -2880 1148
rect -2930 739 -2880 751
rect -2764 1148 -2714 1160
rect -2764 751 -2758 1148
rect -2720 751 -2714 1148
rect -2764 739 -2714 751
rect -2598 1148 -2548 1160
rect -2598 751 -2592 1148
rect -2554 751 -2548 1148
rect -2598 739 -2548 751
rect -2432 1148 -2382 1160
rect -2432 751 -2426 1148
rect -2388 751 -2382 1148
rect -2432 739 -2382 751
rect -2266 1148 -2216 1160
rect -2266 751 -2260 1148
rect -2222 751 -2216 1148
rect -2266 739 -2216 751
rect -2100 1148 -2050 1160
rect -2100 751 -2094 1148
rect -2056 751 -2050 1148
rect -2100 739 -2050 751
rect -1934 1148 -1884 1160
rect -1934 751 -1928 1148
rect -1890 751 -1884 1148
rect -1934 739 -1884 751
rect -1768 1148 -1718 1160
rect -1768 751 -1762 1148
rect -1724 751 -1718 1148
rect -1768 739 -1718 751
rect -1602 1148 -1552 1160
rect -1602 751 -1596 1148
rect -1558 751 -1552 1148
rect -1602 739 -1552 751
rect -1436 1148 -1386 1160
rect -1436 751 -1430 1148
rect -1392 751 -1386 1148
rect -1436 739 -1386 751
rect -1270 1148 -1220 1160
rect -1270 751 -1264 1148
rect -1226 751 -1220 1148
rect -1270 739 -1220 751
rect -1104 1148 -1054 1160
rect -1104 751 -1098 1148
rect -1060 751 -1054 1148
rect -1104 739 -1054 751
rect -938 1148 -888 1160
rect -938 751 -932 1148
rect -894 751 -888 1148
rect -938 739 -888 751
rect -772 1148 -722 1160
rect -772 751 -766 1148
rect -728 751 -722 1148
rect -772 739 -722 751
rect -606 1148 -556 1160
rect -606 751 -600 1148
rect -562 751 -556 1148
rect -606 739 -556 751
rect -440 1148 -390 1160
rect -440 751 -434 1148
rect -396 751 -390 1148
rect -440 739 -390 751
rect -274 1148 -224 1160
rect -274 751 -268 1148
rect -230 751 -224 1148
rect -274 739 -224 751
rect -108 1148 -58 1160
rect -108 751 -102 1148
rect -64 751 -58 1148
rect -108 739 -58 751
rect 58 1148 108 1160
rect 58 751 64 1148
rect 102 751 108 1148
rect 58 739 108 751
rect 224 1148 274 1160
rect 224 751 230 1148
rect 268 751 274 1148
rect 224 739 274 751
rect 390 1148 440 1160
rect 390 751 396 1148
rect 434 751 440 1148
rect 390 739 440 751
rect 556 1148 606 1160
rect 556 751 562 1148
rect 600 751 606 1148
rect 556 739 606 751
rect 722 1148 772 1160
rect 722 751 728 1148
rect 766 751 772 1148
rect 722 739 772 751
rect 888 1148 938 1160
rect 888 751 894 1148
rect 932 751 938 1148
rect 888 739 938 751
rect 1054 1148 1104 1160
rect 1054 751 1060 1148
rect 1098 751 1104 1148
rect 1054 739 1104 751
rect 1220 1148 1270 1160
rect 1220 751 1226 1148
rect 1264 751 1270 1148
rect 1220 739 1270 751
rect 1386 1148 1436 1160
rect 1386 751 1392 1148
rect 1430 751 1436 1148
rect 1386 739 1436 751
rect 1552 1148 1602 1160
rect 1552 751 1558 1148
rect 1596 751 1602 1148
rect 1552 739 1602 751
rect 1718 1148 1768 1160
rect 1718 751 1724 1148
rect 1762 751 1768 1148
rect 1718 739 1768 751
rect 1884 1148 1934 1160
rect 1884 751 1890 1148
rect 1928 751 1934 1148
rect 1884 739 1934 751
rect 2050 1148 2100 1160
rect 2050 751 2056 1148
rect 2094 751 2100 1148
rect 2050 739 2100 751
rect 2216 1148 2266 1160
rect 2216 751 2222 1148
rect 2260 751 2266 1148
rect 2216 739 2266 751
rect 2382 1148 2432 1160
rect 2382 751 2388 1148
rect 2426 751 2432 1148
rect 2382 739 2432 751
rect 2548 1148 2598 1160
rect 2548 751 2554 1148
rect 2592 751 2598 1148
rect 2548 739 2598 751
rect 2714 1148 2764 1160
rect 2714 751 2720 1148
rect 2758 751 2764 1148
rect 2714 739 2764 751
rect 2880 1148 2930 1160
rect 2880 751 2886 1148
rect 2924 751 2930 1148
rect 2880 739 2930 751
rect 3046 1148 3096 1160
rect 3046 751 3052 1148
rect 3090 751 3096 1148
rect 3046 739 3096 751
rect 3212 1148 3262 1160
rect 3212 751 3218 1148
rect 3256 751 3262 1148
rect 3212 739 3262 751
rect 3378 1148 3428 1160
rect 3378 751 3384 1148
rect 3422 751 3428 1148
rect 3378 739 3428 751
rect 3544 1148 3594 1160
rect 3544 751 3550 1148
rect 3588 751 3594 1148
rect 3544 739 3594 751
rect 3710 1148 3760 1160
rect 3710 751 3716 1148
rect 3754 751 3760 1148
rect 3710 739 3760 751
rect 3876 1148 3926 1160
rect 3876 751 3882 1148
rect 3920 751 3926 1148
rect 3876 739 3926 751
rect 4042 1148 4092 1160
rect 4042 751 4048 1148
rect 4086 751 4092 1148
rect 4042 739 4092 751
rect 4208 1148 4258 1160
rect 4208 751 4214 1148
rect 4252 751 4258 1148
rect 4208 739 4258 751
rect 4374 1148 4424 1160
rect 4374 751 4380 1148
rect 4418 751 4424 1148
rect 4374 739 4424 751
rect 4540 1148 4590 1160
rect 4540 751 4546 1148
rect 4584 751 4590 1148
rect 4540 739 4590 751
rect 4706 1148 4756 1160
rect 4706 751 4712 1148
rect 4750 751 4756 1148
rect 4706 739 4756 751
rect 4872 1148 4922 1160
rect 4872 751 4878 1148
rect 4916 751 4922 1148
rect 4872 739 4922 751
rect -4922 -751 -4872 -739
rect -4922 -1148 -4916 -751
rect -4878 -1148 -4872 -751
rect -4922 -1160 -4872 -1148
rect -4756 -751 -4706 -739
rect -4756 -1148 -4750 -751
rect -4712 -1148 -4706 -751
rect -4756 -1160 -4706 -1148
rect -4590 -751 -4540 -739
rect -4590 -1148 -4584 -751
rect -4546 -1148 -4540 -751
rect -4590 -1160 -4540 -1148
rect -4424 -751 -4374 -739
rect -4424 -1148 -4418 -751
rect -4380 -1148 -4374 -751
rect -4424 -1160 -4374 -1148
rect -4258 -751 -4208 -739
rect -4258 -1148 -4252 -751
rect -4214 -1148 -4208 -751
rect -4258 -1160 -4208 -1148
rect -4092 -751 -4042 -739
rect -4092 -1148 -4086 -751
rect -4048 -1148 -4042 -751
rect -4092 -1160 -4042 -1148
rect -3926 -751 -3876 -739
rect -3926 -1148 -3920 -751
rect -3882 -1148 -3876 -751
rect -3926 -1160 -3876 -1148
rect -3760 -751 -3710 -739
rect -3760 -1148 -3754 -751
rect -3716 -1148 -3710 -751
rect -3760 -1160 -3710 -1148
rect -3594 -751 -3544 -739
rect -3594 -1148 -3588 -751
rect -3550 -1148 -3544 -751
rect -3594 -1160 -3544 -1148
rect -3428 -751 -3378 -739
rect -3428 -1148 -3422 -751
rect -3384 -1148 -3378 -751
rect -3428 -1160 -3378 -1148
rect -3262 -751 -3212 -739
rect -3262 -1148 -3256 -751
rect -3218 -1148 -3212 -751
rect -3262 -1160 -3212 -1148
rect -3096 -751 -3046 -739
rect -3096 -1148 -3090 -751
rect -3052 -1148 -3046 -751
rect -3096 -1160 -3046 -1148
rect -2930 -751 -2880 -739
rect -2930 -1148 -2924 -751
rect -2886 -1148 -2880 -751
rect -2930 -1160 -2880 -1148
rect -2764 -751 -2714 -739
rect -2764 -1148 -2758 -751
rect -2720 -1148 -2714 -751
rect -2764 -1160 -2714 -1148
rect -2598 -751 -2548 -739
rect -2598 -1148 -2592 -751
rect -2554 -1148 -2548 -751
rect -2598 -1160 -2548 -1148
rect -2432 -751 -2382 -739
rect -2432 -1148 -2426 -751
rect -2388 -1148 -2382 -751
rect -2432 -1160 -2382 -1148
rect -2266 -751 -2216 -739
rect -2266 -1148 -2260 -751
rect -2222 -1148 -2216 -751
rect -2266 -1160 -2216 -1148
rect -2100 -751 -2050 -739
rect -2100 -1148 -2094 -751
rect -2056 -1148 -2050 -751
rect -2100 -1160 -2050 -1148
rect -1934 -751 -1884 -739
rect -1934 -1148 -1928 -751
rect -1890 -1148 -1884 -751
rect -1934 -1160 -1884 -1148
rect -1768 -751 -1718 -739
rect -1768 -1148 -1762 -751
rect -1724 -1148 -1718 -751
rect -1768 -1160 -1718 -1148
rect -1602 -751 -1552 -739
rect -1602 -1148 -1596 -751
rect -1558 -1148 -1552 -751
rect -1602 -1160 -1552 -1148
rect -1436 -751 -1386 -739
rect -1436 -1148 -1430 -751
rect -1392 -1148 -1386 -751
rect -1436 -1160 -1386 -1148
rect -1270 -751 -1220 -739
rect -1270 -1148 -1264 -751
rect -1226 -1148 -1220 -751
rect -1270 -1160 -1220 -1148
rect -1104 -751 -1054 -739
rect -1104 -1148 -1098 -751
rect -1060 -1148 -1054 -751
rect -1104 -1160 -1054 -1148
rect -938 -751 -888 -739
rect -938 -1148 -932 -751
rect -894 -1148 -888 -751
rect -938 -1160 -888 -1148
rect -772 -751 -722 -739
rect -772 -1148 -766 -751
rect -728 -1148 -722 -751
rect -772 -1160 -722 -1148
rect -606 -751 -556 -739
rect -606 -1148 -600 -751
rect -562 -1148 -556 -751
rect -606 -1160 -556 -1148
rect -440 -751 -390 -739
rect -440 -1148 -434 -751
rect -396 -1148 -390 -751
rect -440 -1160 -390 -1148
rect -274 -751 -224 -739
rect -274 -1148 -268 -751
rect -230 -1148 -224 -751
rect -274 -1160 -224 -1148
rect -108 -751 -58 -739
rect -108 -1148 -102 -751
rect -64 -1148 -58 -751
rect -108 -1160 -58 -1148
rect 58 -751 108 -739
rect 58 -1148 64 -751
rect 102 -1148 108 -751
rect 58 -1160 108 -1148
rect 224 -751 274 -739
rect 224 -1148 230 -751
rect 268 -1148 274 -751
rect 224 -1160 274 -1148
rect 390 -751 440 -739
rect 390 -1148 396 -751
rect 434 -1148 440 -751
rect 390 -1160 440 -1148
rect 556 -751 606 -739
rect 556 -1148 562 -751
rect 600 -1148 606 -751
rect 556 -1160 606 -1148
rect 722 -751 772 -739
rect 722 -1148 728 -751
rect 766 -1148 772 -751
rect 722 -1160 772 -1148
rect 888 -751 938 -739
rect 888 -1148 894 -751
rect 932 -1148 938 -751
rect 888 -1160 938 -1148
rect 1054 -751 1104 -739
rect 1054 -1148 1060 -751
rect 1098 -1148 1104 -751
rect 1054 -1160 1104 -1148
rect 1220 -751 1270 -739
rect 1220 -1148 1226 -751
rect 1264 -1148 1270 -751
rect 1220 -1160 1270 -1148
rect 1386 -751 1436 -739
rect 1386 -1148 1392 -751
rect 1430 -1148 1436 -751
rect 1386 -1160 1436 -1148
rect 1552 -751 1602 -739
rect 1552 -1148 1558 -751
rect 1596 -1148 1602 -751
rect 1552 -1160 1602 -1148
rect 1718 -751 1768 -739
rect 1718 -1148 1724 -751
rect 1762 -1148 1768 -751
rect 1718 -1160 1768 -1148
rect 1884 -751 1934 -739
rect 1884 -1148 1890 -751
rect 1928 -1148 1934 -751
rect 1884 -1160 1934 -1148
rect 2050 -751 2100 -739
rect 2050 -1148 2056 -751
rect 2094 -1148 2100 -751
rect 2050 -1160 2100 -1148
rect 2216 -751 2266 -739
rect 2216 -1148 2222 -751
rect 2260 -1148 2266 -751
rect 2216 -1160 2266 -1148
rect 2382 -751 2432 -739
rect 2382 -1148 2388 -751
rect 2426 -1148 2432 -751
rect 2382 -1160 2432 -1148
rect 2548 -751 2598 -739
rect 2548 -1148 2554 -751
rect 2592 -1148 2598 -751
rect 2548 -1160 2598 -1148
rect 2714 -751 2764 -739
rect 2714 -1148 2720 -751
rect 2758 -1148 2764 -751
rect 2714 -1160 2764 -1148
rect 2880 -751 2930 -739
rect 2880 -1148 2886 -751
rect 2924 -1148 2930 -751
rect 2880 -1160 2930 -1148
rect 3046 -751 3096 -739
rect 3046 -1148 3052 -751
rect 3090 -1148 3096 -751
rect 3046 -1160 3096 -1148
rect 3212 -751 3262 -739
rect 3212 -1148 3218 -751
rect 3256 -1148 3262 -751
rect 3212 -1160 3262 -1148
rect 3378 -751 3428 -739
rect 3378 -1148 3384 -751
rect 3422 -1148 3428 -751
rect 3378 -1160 3428 -1148
rect 3544 -751 3594 -739
rect 3544 -1148 3550 -751
rect 3588 -1148 3594 -751
rect 3544 -1160 3594 -1148
rect 3710 -751 3760 -739
rect 3710 -1148 3716 -751
rect 3754 -1148 3760 -751
rect 3710 -1160 3760 -1148
rect 3876 -751 3926 -739
rect 3876 -1148 3882 -751
rect 3920 -1148 3926 -751
rect 3876 -1160 3926 -1148
rect 4042 -751 4092 -739
rect 4042 -1148 4048 -751
rect 4086 -1148 4092 -751
rect 4042 -1160 4092 -1148
rect 4208 -751 4258 -739
rect 4208 -1148 4214 -751
rect 4252 -1148 4258 -751
rect 4208 -1160 4258 -1148
rect 4374 -751 4424 -739
rect 4374 -1148 4380 -751
rect 4418 -1148 4424 -751
rect 4374 -1160 4424 -1148
rect 4540 -751 4590 -739
rect 4540 -1148 4546 -751
rect 4584 -1148 4590 -751
rect 4540 -1160 4590 -1148
rect 4706 -751 4756 -739
rect 4706 -1148 4712 -751
rect 4750 -1148 4756 -751
rect 4706 -1160 4756 -1148
rect 4872 -751 4922 -739
rect 4872 -1148 4878 -751
rect 4916 -1148 4922 -751
rect 4872 -1160 4922 -1148
<< properties >>
string FIXED_BBOX -5045 -1279 5045 1279
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 7.5 m 1 nx 60 wmin 0.350 lmin 0.50 rho 2000 val 43.932k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
