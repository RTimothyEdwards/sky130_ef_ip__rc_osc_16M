magic
tech sky130A
magscale 1 2
timestamp 1699295625
<< error_s >>
rect 878 76 2736 144
rect 878 -2464 958 76
rect 2418 -836 2736 76
rect 2450 -2258 2736 -836
rect 1164 -2464 2736 -2258
rect 878 -2544 2736 -2464
<< dnwell >>
rect 958 -2464 2656 64
<< nwell >>
rect 958 -148 2418 76
rect 958 -1494 1192 -148
rect 958 -2464 1164 -1494
<< pwell >>
rect -364 -2102 58 -1782
rect 1164 -2454 2458 -1526
<< psubdiff >>
rect -172 -2072 -148 -1978
rect 18 -2072 42 -1978
<< mvpsubdiff >>
rect 1264 -2412 1288 -2316
rect 2394 -2412 2418 -2316
<< psubdiffcont >>
rect -148 -2072 18 -1978
<< mvpsubdiffcont >>
rect 1288 -2412 2394 -2316
<< locali >>
rect 1176 -152 2424 -138
rect 1176 -368 1194 -152
rect 1280 -262 1736 -152
rect 1280 -368 1302 -262
rect -238 -528 -80 -520
rect -238 -612 -220 -528
rect -332 -674 -220 -612
rect -90 -612 -80 -528
rect -90 -674 66 -612
rect -332 -714 66 -674
rect -2 -1180 66 -714
rect 1176 -728 1302 -368
rect 1714 -514 1736 -262
rect 1864 -262 2320 -152
rect 1864 -514 1894 -262
rect 1714 -728 1894 -514
rect 2298 -390 2320 -262
rect 2406 -390 2424 -152
rect 2298 -728 2424 -390
rect 1176 -914 2424 -728
rect -2 -1708 64 -1260
rect 1176 -1380 1302 -914
rect 1714 -1380 1894 -914
rect 2298 -1380 2424 -914
rect 1176 -1488 2424 -1380
rect -334 -1796 64 -1708
rect -334 -1810 -190 -1796
rect -236 -1918 -190 -1810
rect -52 -1810 64 -1796
rect 1184 -1644 2426 -1538
rect -52 -1918 34 -1810
rect -236 -1978 34 -1918
rect -236 -2072 -148 -1978
rect 18 -2072 34 -1978
rect 1184 -2070 1310 -1644
rect 1698 -1980 1914 -1644
rect 1698 -2070 1708 -1980
rect 1184 -2148 1708 -2070
rect 1184 -2212 1356 -2148
rect 1612 -2198 1708 -2148
rect 1904 -2070 1914 -1980
rect 2300 -2070 2426 -1644
rect 1904 -2146 2426 -2070
rect 1904 -2198 1992 -2146
rect 1612 -2210 1992 -2198
rect 2248 -2210 2426 -2146
rect 1612 -2212 2426 -2210
rect 1184 -2236 2426 -2212
rect 1272 -2412 1288 -2316
rect 2394 -2412 2410 -2316
<< viali >>
rect 1194 -368 1280 -152
rect -220 -674 -90 -528
rect 1736 -514 1864 -152
rect 2320 -390 2406 -152
rect -190 -1918 -52 -1796
rect 1356 -2212 1612 -2148
rect 1708 -2198 1904 -1980
rect 1992 -2210 2248 -2146
<< metal1 >>
rect 1174 -152 2426 64
rect 1174 -368 1194 -152
rect 1280 -263 1736 -152
rect 1280 -368 1300 -263
rect 1174 -382 1300 -368
rect -422 -528 56 -520
rect -422 -674 -220 -528
rect -90 -674 56 -528
rect -422 -720 56 -674
rect -254 -996 -208 -720
rect -422 -1166 -222 -1104
rect -186 -1166 -138 -1034
rect -422 -1240 -218 -1166
rect -138 -1240 -128 -1166
rect -422 -1304 -222 -1240
rect -186 -1406 -138 -1240
rect -264 -1714 -218 -1432
rect -96 -1488 -54 -790
rect 1336 -1198 1402 -446
rect 1468 -662 1520 -366
rect 1618 -444 1736 -263
rect 1554 -514 1736 -444
rect 1864 -263 2320 -152
rect 1864 -444 1996 -263
rect 1864 -514 2048 -444
rect 1554 -530 2048 -514
rect 1468 -714 1644 -662
rect 1592 -880 1644 -714
rect 1910 -722 1920 -656
rect 2018 -664 2028 -656
rect 2086 -664 2138 -368
rect 2300 -390 2320 -263
rect 2406 -390 2426 -152
rect 2300 -412 2426 -390
rect 2018 -716 2138 -664
rect 2018 -722 2028 -716
rect 1580 -946 1590 -880
rect 1688 -946 1698 -880
rect 1442 -1076 1452 -1010
rect 1550 -1076 1560 -1010
rect 1482 -1274 1524 -1076
rect 1592 -1230 1644 -946
rect 1962 -1012 2014 -722
rect 1910 -1078 1920 -1012
rect 2018 -1078 2028 -1012
rect 1582 -1296 1592 -1230
rect 1690 -1296 1700 -1230
rect 1408 -1422 1418 -1356
rect 1516 -1422 1526 -1356
rect -96 -1554 -64 -1488
rect 34 -1554 44 -1488
rect -96 -1560 -54 -1554
rect -264 -1726 -216 -1714
rect -396 -1796 52 -1726
rect 1476 -1736 1516 -1422
rect 1456 -1738 1516 -1736
rect -396 -1918 -190 -1796
rect -52 -1918 52 -1796
rect -396 -1926 52 -1918
rect 1336 -2046 1420 -1814
rect 1476 -1962 1516 -1738
rect 1592 -1902 1644 -1296
rect 1962 -1906 2014 -1078
rect 2082 -1230 2124 -1012
rect 2204 -1198 2270 -446
rect 2450 -648 2650 -522
rect 2310 -714 2320 -648
rect 2418 -714 2650 -648
rect 2450 -722 2650 -714
rect 2456 -878 2656 -870
rect 2310 -944 2320 -878
rect 2418 -944 2656 -878
rect 2456 -1070 2656 -944
rect 2052 -1296 2062 -1230
rect 2160 -1296 2170 -1230
rect 2054 -1554 2064 -1488
rect 2162 -1498 2172 -1488
rect 2456 -1498 2656 -1408
rect 2162 -1546 2656 -1498
rect 2162 -1554 2172 -1546
rect 2088 -1964 2128 -1554
rect 2456 -1608 2656 -1546
rect 1652 -1980 1962 -1972
rect 1652 -2046 1708 -1980
rect 1336 -2148 1708 -2046
rect 1336 -2212 1356 -2148
rect 1612 -2198 1708 -2148
rect 1904 -2046 1962 -1980
rect 2184 -2046 2268 -1812
rect 1904 -2146 2268 -2046
rect 1904 -2198 1992 -2146
rect 1612 -2210 1992 -2198
rect 2248 -2210 2268 -2146
rect 1612 -2212 2268 -2210
rect 1336 -2264 2268 -2212
rect 1165 -2464 2653 -2264
<< via1 >>
rect -218 -1240 -138 -1166
rect 1920 -722 2018 -656
rect 1590 -946 1688 -880
rect 1452 -1076 1550 -1010
rect 1920 -1078 2018 -1012
rect 1592 -1296 1690 -1230
rect 1418 -1422 1516 -1356
rect -64 -1554 34 -1488
rect 2320 -714 2418 -648
rect 2320 -944 2418 -878
rect 2062 -1296 2160 -1230
rect 2064 -1554 2162 -1488
<< metal2 >>
rect 1920 -656 2018 -646
rect 2320 -648 2418 -638
rect 2018 -710 2320 -656
rect 1920 -732 2018 -722
rect 2320 -724 2418 -714
rect 1590 -880 1688 -870
rect 2320 -878 2418 -868
rect 1688 -942 2320 -886
rect 1590 -956 1688 -946
rect 2320 -954 2418 -944
rect 1452 -1010 1550 -1000
rect 1920 -1012 2018 -1002
rect 1550 -1072 1920 -1018
rect 1452 -1086 1550 -1076
rect 2018 -1072 2032 -1018
rect 1920 -1088 2018 -1078
rect -218 -1166 -138 -1156
rect -138 -1231 50 -1177
rect -218 -1250 -138 -1240
rect -4 -1364 50 -1231
rect 1592 -1230 1690 -1220
rect 1572 -1286 1592 -1232
rect 2062 -1230 2160 -1220
rect 1690 -1286 2062 -1232
rect 1592 -1306 1690 -1296
rect 2062 -1306 2160 -1296
rect 1418 -1356 1516 -1346
rect -4 -1418 1418 -1364
rect 1418 -1432 1516 -1422
rect -64 -1488 34 -1478
rect 2064 -1488 2162 -1478
rect 34 -1548 2064 -1494
rect -64 -1564 34 -1554
rect 2064 -1564 2162 -1554
use sky130_fd_pr__pfet_01v8_LGS3BL  XM7 paramcells
timestamp 1699295625
transform 1 0 -153 0 1 -932
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_64Z3AY  XM8 paramcells
timestamp 1699295625
transform 1 0 -153 0 1 -1503
box -211 -279 211 279
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM15 paramcells
timestamp 1699295625
transform 1 0 1500 0 1 -1155
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM16
timestamp 1699295625
transform 1 0 1494 0 1 -487
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM17 paramcells
timestamp 1699295625
transform 1 0 1502 0 1 -1858
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM18
timestamp 1699295625
transform 1 0 2108 0 1 -1856
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM19
timestamp 1699295625
transform 1 0 2110 0 1 -487
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM20
timestamp 1699295625
transform 1 0 2110 0 1 -1157
box -308 -339 308 339
<< labels >>
flabel metal1 2450 -722 2650 -522 0 FreeSans 256 0 0 0 out_h
port 1 nsew
flabel metal1 2456 -1070 2656 -870 0 FreeSans 256 0 0 0 outb_h
port 3 nsew
flabel metal1 2456 -1608 2656 -1408 0 FreeSans 256 0 0 0 inb_l
port 7 nsew
flabel metal1 -422 -1304 -222 -1104 0 FreeSans 256 0 0 0 in_l
port 4 nsew
flabel metal1 -396 -1926 -196 -1726 0 FreeSans 256 0 0 0 dvss
port 5 nsew
flabel metal1 -422 -720 -222 -520 0 FreeSans 256 0 0 0 dvdd
port 0 nsew
flabel metal1 2453 -2464 2653 -2264 0 FreeSans 256 0 0 0 avss
port 6 nsew
flabel metal1 2226 -136 2426 64 0 FreeSans 256 0 0 0 avdd
port 2 nsew
<< end >>
