* NGSPICE file created from sky130_ef_ip__rc_osc_16M.ext - technology: sky130A

** x1 ena vdd1v8 vdd3v3 GND GND dout sky130_ef_ip__rc_osc_16M

.subckt sky130_ef_ip__rc_osc_16M ena dvdd avdd dvss avss dout
X0 a_1178_9068# a_1344_7168# avss.t101 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X1 avdd.t19 a_1538_5653.t0 a_1538_5653.t1 avdd.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X2 a_6490_9068# a_6656_7168# avss.t15 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X3 a_7672_3118# a_7506_1218# avss.t8 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X4 a_2360_3118# a_2194_1218# avss.t82 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X5 a_3502_9068# a_3336_7168# avss.t66 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X6 a_5162_9068# a_4996_7168# avss.t14 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X7 a_7008_3118# a_6842_1218# avss.t57 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X8 a_8814_9068# a_8648_7168# avss.t56 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X9 a_2692_3118# a_2858_1218# avss.t55 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X10 avss.t103 ena.t0 rc_osc_level_shifter_0.outb_h.t1 avss.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X11 a_9664_3118# a_9830_1218# avss.t79 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X12 a_9996_3118# a_10162_1218# avss.t76 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X13 a_7154_9068# a_7320_7168# avss.t40 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X14 a_1364_3118# a_1198_1218# avss.t7 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X15 dvdd.t7 ena.t1 rc_osc_level_shifter_0.inb_l dvdd.t6 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X16 a_6676_3118# a_6510_1218# avss.t75 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X17 a_6444_4786# a_2982_4700.t2 avss.t100 avss.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X18 a_4166_9068# a_4000_7168# avss.t78 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X19 a_4194_4788# a_3638_4788# a_4036_4788# avss.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X20 a_2506_9068# a_2340_7168# avss.t49 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X21 a_9478_9068# a_9312_7168# avss.t77 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X22 a_7818_9068# a_7652_7168# avss.t32 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X23 a_5016_3118# a_5182_1218# avss.t31 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X24 a_8668_3118# a_8834_1218# avss.t38 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X25 a_3356_3118# a_3522_1218# avss.t37 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X26 avdd.t15 a_1538_5653.t10 a_1538_5653.t11 avdd.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X27 a_846_9068# a_1012_7168# avss.t71 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X28 a_6158_9068# a_6324_7168# avss.t13 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X29 a_7340_3118# a_7174_1218# avss.t65 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X30 a_10142_9068# a_10308_7168# avss.t25 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X31 avdd.t16 a_1538_5653.t14 a_4854_5653# avdd.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X32 avdd.t18 a_1538_5653.t8 a_1538_5653.t9 avdd.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X33 a_9332_3118# a_9498_1218# avss.t114 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X34 a_4020_3118# a_4186_1218# avss.t112 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X35 a_2360_3118# a_2526_1218# avss.t29 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X36 a_5826_9068# a_5992_7168# avss.t45 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X37 a_7672_3118# a_7838_1218# avss.t36 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X38 a_5162_9068# a_5328_7168# avss.t136 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X39 dvss.t6 ena.t2 rc_osc_level_shifter_0.inb_l dvss.t5 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X40 avdd.t13 a_1538_5653.t15 a_5470_5653# avdd.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X41 a_1032_3118# a_866_1218# avss.t64 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X42 a_6344_3118# a_6178_1218# avss.t48 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X43 a_6602_4786# ena.t3 a_6444_4786# avss.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X44 a_1538_5653.t7 a_1538_5653.t6 avdd.t11 avdd.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X45 a_9146_9068# a_8980_7168# avss.t63 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X46 a_10308_7168# a_10162_1218# avss.t135 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X47 a_4830_9068# a_4996_7168# avss.t27 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X48 a_8336_3118# a_8502_1218# avss.t85 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X49 a_5348_3118# a_5182_1218# avss.t24 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X50 a_1842_9068# a_1676_7168# avss.t54 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X51 avdd.t28 rc_osc_level_shifter_0.out_h.t2 a_1538_5653.t12 avdd.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X52 a_9000_3118# a_9166_1218# avss.t81 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X53 a_5494_9068# a_5660_7168# avss.t80 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X54 a_7340_3118# a_7506_1218# avss.t122 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X55 a_4750_4788# a_4194_4788# a_4854_5653# avdd.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X56 a_1414_4786.t3 rc_osc_level_shifter_0.outb_h.t2 avss.t47 avss.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X57 avdd.t10 a_1538_5653.t4 a_1538_5653.t5 avdd.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X58 a_6012_3118# a_5846_1218# avss.t28 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X59 a_8366_5327# rc_osc_level_shifter_0.out_h.t3 rc_osc_level_shifter_0.outb_h.t0 avdd.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X60 a_1696_3118# a_1862_1218# avss.t113 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X61 a_1414_4786.t2 rc_osc_level_shifter_0.out_h.t4 a_514_7168.t1 avss.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X62 a_700_3118# a_534_1218# avss.t23 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X63 a_2982_4700.t1 a_4750_4788# a_5470_5653# avdd.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X64 a_4498_9068# a_4664_7168# avss.t53 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X65 a_9810_9068# a_9976_7168# avss.t98 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X66 avdd.t4 a_1538_5653.t16 a_3622_5653# avdd.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X67 a_1538_5653.t3 a_1538_5653.t2 avdd.t8 avdd.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X68 a_5680_3118# a_5514_1218# avss.t39 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X69 a_3170_9068# a_3004_7168# avss.t22 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X70 a_5016_3118# a_4850_1218# avss.t68 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X71 a_1510_9068# a_1344_7168# avss.t130 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X72 a_6822_9068# a_6656_7168# avss.t111 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X73 a_8482_9068# a_8316_7168# avss.t117 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X74 avdd.t6 a_1538_5653.t17 a_3006_5653# avdd.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X75 dout.t0 a_6602_4786# dvss.t1 dvss.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
X76 avdd.t2 a_1538_5653.t18 a_4238_5653# avdd.t1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X77 a_3502_9068# a_3668_7168# avss.t26 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X78 rc_osc_level_shifter_0.out_h.t1 rc_osc_level_shifter_0.outb_h.t3 a_7598_4659# avdd.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X79 rc_osc_level_shifter_0.out_h.t0 rc_osc_level_shifter_0.inb_l avss.t52 avss.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X80 a_9996_3118# a_9830_1218# avss.t62 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X81 a_4684_3118# a_4518_1218# avss.t86 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X82 a_2174_9068# a_2008_7168# avss.t17 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X83 a_7486_9068# a_7320_7168# avss.t30 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X84 dout.t1 rc_osc_level_shifter_0.inb_l a_10681_5200# dvdd.t2 sky130_fd_pr__pfet_01v8 ad=0.465 pd=3.62 as=0.2475 ps=1.83 w=1.5 l=0.15
X85 a_5826_9068# a_5660_7168# avss.t74 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X86 a_3024_3118# a_3190_1218# avss.t134 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X87 a_1364_3118# a_1530_1218# avss.t84 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X88 a_6676_3118# a_6842_1218# avss.t44 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X89 a_4166_9068# a_4332_7168# avss.t21 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X90 a_9478_9068# a_9644_7168# avss.t73 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X91 a_3688_3118# a_3522_1218# avss.t124 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X92 a_514_9068# a_680_7168# avss.t20 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X93 a_1178_9068# a_1012_7168# avss.t19 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X94 a_5148_4788# a_1414_4786.t4 avss.t97 avss.t96 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X95 a_8150_9068# a_7984_7168# avss.t129 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X96 a_2028_3118# a_2194_1218# avss.t70 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X97 a_5680_3118# a_5846_1218# avss.t139 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X98 a_6602_4786# a_2982_4700.t3 dvdd.t3 avdd.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.5
X99 a_3638_4788# a_3082_4788# a_3622_5653# avdd.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X100 a_3480_4788# a_1414_4786.t5 avss.t95 avss.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X101 a_3170_9068# a_3336_7168# avss.t141 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X102 a_8482_9068# a_8648_7168# avss.t69 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X103 a_3082_4788# a_2982_4700.t4 a_3006_5653# avdd.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X104 a_4352_3118# a_4186_1218# avss.t138 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X105 a_9664_3118# a_9498_1218# avss.t131 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X106 dvss.t4 ena.t4 sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
X107 a_4194_4788# a_3638_4788# a_4238_5653# avdd.t1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X108 a_7154_9068# a_6988_7168# avss.t140 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X109 a_1032_3118# a_1198_1218# avss.t128 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X110 a_8004_3118# a_8170_1218# avss.t12 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X111 avdd.t29 rc_osc_level_shifter_0.out_h.t5 a_7598_4659# avdd.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X112 a_6344_3118# a_6510_1218# avss.t127 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X113 a_3834_9068# a_4000_7168# avss.t120 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X114 a_9146_9068# a_9312_7168# avss.t72 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X115 a_3356_3118# a_3190_1218# avss.t133 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X116 a_8668_3118# a_8502_1218# avss.t137 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X117 dvss.t3 rc_osc_level_shifter_0.inb_l dout.t2 dvss.t2 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X118 a_6158_9068# a_5992_7168# avss.t67 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X119 a_2982_4700.t0 a_4750_4788# a_5148_4788# avss.t96 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X120 a_4592_4788# a_1414_4786.t6 avss.t92 avss.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X121 a_7008_3118# a_7174_1218# avss.t121 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X122 a_5348_3118# a_5514_1218# avss.t83 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X123 a_846_9068# a_680_7168# avss.t123 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X124 a_8814_9068# a_8980_7168# avss.t11 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X125 avdd.t22 a_3004_7168# avss.t61 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X126 a_8150_9068# a_8316_7168# avss.t132 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X127 a_2526_4188# a_1414_4786.t7 avss.t91 avss.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X128 a_3638_4788# a_3082_4788# a_3480_4788# avss.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X129 a_4020_3118# a_3854_1218# avss.t110 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X130 a_2924_4788# a_1414_4786.t8 avss.t89 avss.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X131 a_9332_3118# a_9166_1218# avss.t5 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X132 a_6012_3118# a_6178_1218# avss.t4 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X133 a_2506_9068# a_2672_7168# avss.t109 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X134 a_7818_9068# a_7984_7168# avss.t119 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X135 a_4352_3118# a_4518_1218# avss.t118 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X136 dvdd.t5 ena.t5 a_6602_4786# dvdd.t4 sky130_fd_pr__pfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X137 a_1842_9068# a_2008_7168# avss.t3 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X138 a_700_3118# a_866_1218# avss.t2 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X139 a_6490_9068# a_6324_7168# avss.t108 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X140 a_8336_3118# a_8170_1218# avss.t93 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X141 a_3024_3118# a_2858_1218# avss.t10 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X142 a_4830_9068# a_4664_7168# avss.t43 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X143 a_1510_9068# a_1676_7168# avss.t1 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X144 a_514_9068# a_514_7168.t0 avss.t0 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X145 a_6822_9068# a_6988_7168# avss.t116 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X146 a_4750_4788# a_4194_4788# a_4592_4788# avss.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X147 a_2692_3118# a_2526_1218# avss.t106 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X148 a_2028_3118# a_1862_1218# avss.t105 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X149 a_5494_9068# a_5328_7168# avss.t104 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X150 a_9000_3118# a_8834_1218# avss.t60 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X151 a_2526_4188# rc_osc_level_shifter_0.out_h.t6 a_1538_5653.t13 avss.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X152 a_3834_9068# a_3668_7168# avss.t35 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X153 a_1414_4786.t1 a_1414_4786.t0 avss.t99 avss.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X154 a_3082_4788# a_2982_4700.t5 a_2924_4788# avss.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X155 a_4684_3118# a_4850_1218# avss.t9 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X156 a_2174_9068# a_2340_7168# avss.t34 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X157 a_7486_9068# a_7652_7168# avss.t16 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X158 a_1696_3118# a_1530_1218# avss.t107 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X159 avdd.t21 a_534_1218# avss.t59 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X160 a_4036_4788# a_1414_4786.t9 avss.t115 avss.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X161 a_8366_5327# rc_osc_level_shifter_0.outb_h.t4 avdd.t25 avdd.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X162 avdd.t20 a_2672_7168# avss.t42 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X163 a_4498_9068# a_4332_7168# avss.t58 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X164 a_8004_3118# a_7838_1218# avss.t18 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X165 a_9810_9068# a_9644_7168# avss.t41 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X166 a_3688_3118# a_3854_1218# avss.t126 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X167 a_10681_5200# a_6602_4786# dvdd.t1 dvdd.t0 sky130_fd_pr__pfet_01v8 ad=0.2475 pd=1.83 as=0.465 ps=3.62 w=1.5 l=0.15
X168 a_10142_9068# a_9976_7168# avss.t125 sky130_fd_pr__res_xhigh_po_0p35 l=7.5
R0 avss.n200 avss.n3 36543.5
R1 avss.n290 avss.n3 36543.5
R2 avss.n200 avss.n4 36543.5
R3 avss.n290 avss.n4 36543.5
R4 avss.n287 avss.n5 36543.5
R5 avss.n287 avss.n6 36543.5
R6 avss.n12 avss.n6 36543.5
R7 avss.n12 avss.n5 36543.5
R8 avss.t51 avss.n264 10971.7
R9 avss.t102 avss.n14 7496.3
R10 avss.n289 avss.n288 5872.44
R11 avss.t102 avss.n11 1380.27
R12 avss.n279 avss.n15 1379.81
R13 avss.n279 avss.n16 1379.81
R14 avss.n266 avss.n16 1379.81
R15 avss.n217 avss.n83 1379.81
R16 avss.n216 avss.n83 1379.81
R17 avss.n216 avss.n82 1379.81
R18 avss.n217 avss.n82 1379.81
R19 avss.n222 avss.n76 1379.81
R20 avss.n223 avss.n76 1379.81
R21 avss.n223 avss.n75 1379.81
R22 avss.n222 avss.n75 1379.81
R23 avss.n180 avss.n151 1379.81
R24 avss.n179 avss.n151 1379.81
R25 avss.n179 avss.n150 1379.81
R26 avss.n180 avss.n150 1379.81
R27 avss.n185 avss.n145 1379.81
R28 avss.n145 avss.n140 1379.81
R29 avss.n144 avss.n140 1379.81
R30 avss.n185 avss.n144 1379.81
R31 avss.n234 avss.n60 1379.81
R32 avss.n233 avss.n60 1379.81
R33 avss.n233 avss.n59 1379.81
R34 avss.n234 avss.n59 1379.81
R35 avss.n239 avss.n53 1379.81
R36 avss.n240 avss.n53 1379.81
R37 avss.n240 avss.n52 1379.81
R38 avss.n239 avss.n52 1379.81
R39 avss.n121 avss.n100 1379.81
R40 avss.n100 avss.n95 1379.81
R41 avss.n96 avss.n95 1379.81
R42 avss.n121 avss.n96 1379.81
R43 avss.n115 avss.n34 1379.81
R44 avss.n115 avss.n35 1379.81
R45 avss.n253 avss.n35 1379.81
R46 avss.n253 avss.n34 1379.81
R47 avss.n168 avss.n73 1379.81
R48 avss.n168 avss.n77 1379.81
R49 avss.n176 avss.n77 1379.81
R50 avss.n176 avss.n73 1379.81
R51 avss.n175 avss.n152 1379.81
R52 avss.n175 avss.n174 1379.81
R53 avss.n174 avss.n155 1379.81
R54 avss.n155 avss.n152 1379.81
R55 avss.n139 avss.n138 1379.81
R56 avss.n186 avss.n138 1379.81
R57 avss.n186 avss.n137 1379.81
R58 avss.n139 avss.n137 1379.81
R59 avss.n141 avss.n61 1379.81
R60 avss.n141 avss.n62 1379.81
R61 avss.n132 avss.n62 1379.81
R62 avss.n132 avss.n61 1379.81
R63 avss.n129 avss.n49 1379.81
R64 avss.n129 avss.n54 1379.81
R65 avss.n97 avss.n54 1379.81
R66 avss.n97 avss.n49 1379.81
R67 avss.n94 avss.n93 1379.81
R68 avss.n122 avss.n93 1379.81
R69 avss.n122 avss.n92 1379.81
R70 avss.n94 avss.n92 1379.81
R71 avss.n112 avss.n39 1379.81
R72 avss.n112 avss.n104 1379.81
R73 avss.n104 avss.n32 1379.81
R74 avss.n39 avss.n32 1379.81
R75 avss.n255 avss.n25 1379.81
R76 avss.n255 avss.n26 1379.81
R77 avss.n262 avss.n26 1379.81
R78 avss.n262 avss.n25 1379.81
R79 avss.n257 avss.n30 1379.81
R80 avss.n31 avss.n30 1379.81
R81 avss.n31 avss.n24 1379.81
R82 avss.n257 avss.n24 1379.81
R83 avss.n273 avss.n21 1379.81
R84 avss.n275 avss.n20 1379.81
R85 avss.n275 avss.n21 1379.81
R86 avss.n280 avss.n14 1030.34
R87 avss.n281 avss.n11 816.495
R88 avss.n8 avss.n7 712.534
R89 avss.n201 avss.n2 710.625
R90 avss.n286 avss.n7 701.706
R91 avss.n291 avss.n2 691.966
R92 avss.n274 avss.n20 683.336
R93 avss.n266 avss.n265 683.336
R94 avss.n286 avss.n285 627.799
R95 avss.n202 avss.n199 516.365
R96 avss.n284 avss.n8 434.414
R97 avss.n281 avss.n280 349.926
R98 avss.n292 avss.n1 318.509
R99 avss.n285 avss.n284 276.212
R100 avss.t135 avss.t76 267.938
R101 avss.t76 avss.t62 267.938
R102 avss.t62 avss.t79 267.938
R103 avss.t79 avss.t131 267.938
R104 avss.t131 avss.t114 267.938
R105 avss.t114 avss.t5 267.938
R106 avss.t5 avss.t81 267.938
R107 avss.t81 avss.t60 267.938
R108 avss.t60 avss.t38 267.938
R109 avss.t38 avss.t137 267.938
R110 avss.t125 avss.t25 267.546
R111 avss.t98 avss.t125 267.546
R112 avss.t41 avss.t98 267.546
R113 avss.t73 avss.t41 267.546
R114 avss.t77 avss.t73 267.546
R115 avss.t72 avss.t77 267.546
R116 avss.t63 avss.t72 267.546
R117 avss.t11 avss.t63 267.546
R118 avss.t56 avss.t11 267.546
R119 avss.t69 avss.t56 267.546
R120 avss.n200 avss.t135 255.6
R121 avss.t25 avss.n12 255.25
R122 avss.n198 avss.n1 248.393
R123 avss.t137 avss.t85 244.707
R124 avss.t132 avss.t117 244.363
R125 avss.t129 avss.t132 244.363
R126 avss.t119 avss.t129 244.363
R127 avss.t32 avss.t119 244.363
R128 avss.t16 avss.t30 244.363
R129 avss.t30 avss.t40 244.363
R130 avss.t40 avss.t140 244.363
R131 avss.t140 avss.t116 244.363
R132 avss.t116 avss.t111 244.363
R133 avss.t111 avss.t15 244.363
R134 avss.t15 avss.t108 244.363
R135 avss.t108 avss.t13 244.363
R136 avss.t13 avss.t67 244.363
R137 avss.t67 avss.t45 244.363
R138 avss.t74 avss.t80 244.281
R139 avss.t80 avss.t104 244.281
R140 avss.t136 avss.t14 244.281
R141 avss.t14 avss.t27 244.281
R142 avss.t27 avss.t43 244.281
R143 avss.t43 avss.t53 244.281
R144 avss.t53 avss.t58 244.281
R145 avss.t58 avss.t21 244.281
R146 avss.t21 avss.t78 244.281
R147 avss.t78 avss.t120 244.281
R148 avss.t120 avss.t35 244.281
R149 avss.t35 avss.t26 244.281
R150 avss.t26 avss.t66 244.281
R151 avss.t66 avss.t141 244.281
R152 avss.t141 avss.t22 244.281
R153 avss.t22 avss.t61 244.281
R154 avss.t61 avss.t42 244.281
R155 avss.t42 avss.t109 244.281
R156 avss.t109 avss.t49 244.281
R157 avss.t49 avss.t34 244.281
R158 avss.t34 avss.t17 244.281
R159 avss.t17 avss.t3 244.281
R160 avss.t3 avss.t54 244.281
R161 avss.t54 avss.t1 244.281
R162 avss.t1 avss.t130 244.281
R163 avss.t130 avss.t101 244.281
R164 avss.t101 avss.t19 244.281
R165 avss.t19 avss.t71 244.281
R166 avss.t71 avss.t123 244.281
R167 avss.t20 avss.t0 244.281
R168 avss.t51 avss.n14 236.889
R169 avss.n41 avss.t100 235.553
R170 avss.t0 avss.n287 234.507
R171 avss.t85 avss.t93 234.404
R172 avss.t93 avss.t12 234.404
R173 avss.t12 avss.t18 234.404
R174 avss.t18 avss.t36 234.404
R175 avss.t36 avss.t8 234.404
R176 avss.t8 avss.t122 234.404
R177 avss.n213 avss.t47 234.381
R178 avss.n66 avss.t89 234.012
R179 avss.n230 avss.t95 234.012
R180 avss.n50 avss.t115 234.012
R181 avss.n245 avss.t92 234.012
R182 avss.n248 avss.t97 234.012
R183 avss.n228 avss.t91 234.012
R184 avss.n86 avss.t99 233.994
R185 avss.n22 avss.t103 233.939
R186 avss.n88 avss.t52 233.929
R187 avss.t45 avss.t74 225.959
R188 avss.t117 avss.t69 222.579
R189 avss.t122 avss.t65 215.56
R190 avss.t65 avss.t121 169.584
R191 avss.t57 avss.t44 169.584
R192 avss.t127 avss.t48 169.584
R193 avss.n288 avss.t20 169.232
R194 avss.t4 avss.t28 168.529
R195 avss.t28 avss.t139 168.529
R196 avss.t139 avss.t39 168.529
R197 avss.t39 avss.t83 168.529
R198 avss.t31 avss.t68 168.529
R199 avss.t9 avss.t86 168.529
R200 avss.t133 avss.t37 168.529
R201 avss.t134 avss.t10 168.529
R202 avss.t107 avss.t113 168.529
R203 avss.t84 avss.t7 168.529
R204 avss.t64 avss.t2 168.529
R205 avss.t59 avss.t23 168.529
R206 avss.n290 avss.t59 166.969
R207 avss.t87 avss.t75 162.434
R208 avss.t6 avss.t118 149.239
R209 avss.n258 avss.n257 146.25
R210 avss.n257 avss.t87 146.25
R211 avss.n106 avss.n31 146.25
R212 avss.t87 avss.n31 146.25
R213 avss.n260 avss.n25 146.25
R214 avss.t87 avss.n25 146.25
R215 avss.n258 avss.n26 146.25
R216 avss.t87 avss.n26 146.25
R217 avss.n250 avss.n39 146.25
R218 avss.t96 avss.n39 146.25
R219 avss.n109 avss.n104 146.25
R220 avss.n104 avss.t96 146.25
R221 avss.n94 avss.n44 146.25
R222 avss.t6 avss.n94 146.25
R223 avss.n123 avss.n122 146.25
R224 avss.n122 avss.t6 146.25
R225 avss.n241 avss.n49 146.25
R226 avss.t50 avss.n49 146.25
R227 avss.n126 avss.n54 146.25
R228 avss.t50 avss.n54 146.25
R229 avss.n232 avss.n61 146.25
R230 avss.t94 avss.n61 146.25
R231 avss.n190 avss.n62 146.25
R232 avss.t94 avss.n62 146.25
R233 avss.n159 avss.n139 146.25
R234 avss.t88 avss.n139 146.25
R235 avss.n187 avss.n186 146.25
R236 avss.n186 avss.t88 146.25
R237 avss.n152 avss.n68 146.25
R238 avss.t90 avss.n152 146.25
R239 avss.n174 avss.n173 146.25
R240 avss.t90 avss.n174 146.25
R241 avss.n224 avss.n73 146.25
R242 avss.t33 avss.n73 146.25
R243 avss.n170 avss.n77 146.25
R244 avss.t33 avss.n77 146.25
R245 avss.n38 avss.n34 146.25
R246 avss.t96 avss.n34 146.25
R247 avss.n250 avss.n35 146.25
R248 avss.t96 avss.n35 146.25
R249 avss.n121 avss.n120 146.25
R250 avss.t6 avss.n121 146.25
R251 avss.n95 avss.n44 146.25
R252 avss.t6 avss.n95 146.25
R253 avss.n239 avss.n238 146.25
R254 avss.t50 avss.n239 146.25
R255 avss.n241 avss.n240 146.25
R256 avss.n240 avss.t50 146.25
R257 avss.n235 avss.n234 146.25
R258 avss.n234 avss.t94 146.25
R259 avss.n233 avss.n232 146.25
R260 avss.t94 avss.n233 146.25
R261 avss.n185 avss.n184 146.25
R262 avss.t88 avss.n185 146.25
R263 avss.n159 avss.n140 146.25
R264 avss.t88 avss.n140 146.25
R265 avss.n181 avss.n180 146.25
R266 avss.n180 avss.t90 146.25
R267 avss.n179 avss.n68 146.25
R268 avss.t90 avss.n179 146.25
R269 avss.n222 avss.n221 146.25
R270 avss.t33 avss.n222 146.25
R271 avss.n224 avss.n223 146.25
R272 avss.n223 avss.t33 146.25
R273 avss.n218 avss.n217 146.25
R274 avss.n217 avss.t46 146.25
R275 avss.n216 avss.n215 146.25
R276 avss.t46 avss.n216 146.25
R277 avss.n18 avss.n16 146.25
R278 avss.t51 avss.n16 146.25
R279 avss.n269 avss.n15 146.25
R280 avss.n276 avss.n275 146.25
R281 avss.n275 avss.t102 146.25
R282 avss.n273 avss.n272 146.25
R283 avss.t33 avss.t105 145.179
R284 avss.t88 avss.t55 141.118
R285 avss.n98 avss.t112 138.071
R286 avss.t94 avss.t124 137.056
R287 avss.t82 avss.n178 134.011
R288 avss.n14 avss.t32 133.958
R289 avss.t46 avss.t128 132.995
R290 avss.n114 avss.n113 131.981
R291 avss.n143 avss.n142 131.981
R292 avss.n167 avss.n166 131.981
R293 avss.n154 avss.t29 129.95
R294 avss.t96 avss.t24 128.935
R295 avss.n256 avss.t4 128.472
R296 avss.n130 avss.t110 125.888
R297 avss.t104 avss.n13 122.141
R298 avss.n13 avss.t136 122.141
R299 avss.n105 avss.n24 117.207
R300 avss.n263 avss.n24 117.001
R301 avss.n30 avss.n28 117.001
R302 avss.n256 avss.n30 117.001
R303 avss.n262 avss.n261 117.001
R304 avss.n263 avss.n262 117.001
R305 avss.n255 avss.n29 117.001
R306 avss.n256 avss.n255 117.001
R307 avss.n36 avss.n32 117.001
R308 avss.n254 avss.n32 117.001
R309 avss.n112 avss.n111 117.001
R310 avss.n114 avss.n112 117.001
R311 avss.n101 avss.n92 117.001
R312 avss.n113 avss.n92 117.001
R313 avss.n93 avss.n46 117.001
R314 avss.n99 avss.n93 117.001
R315 avss.n97 avss.n48 117.001
R316 avss.n98 avss.n97 117.001
R317 avss.n129 avss.n128 117.001
R318 avss.n130 avss.n129 117.001
R319 avss.n133 avss.n132 117.001
R320 avss.n132 avss.n131 117.001
R321 avss.n141 avss.n134 117.001
R322 avss.n142 avss.n141 117.001
R323 avss.n137 avss.n135 117.001
R324 avss.n143 avss.n137 117.001
R325 avss.n156 avss.n138 117.001
R326 avss.n153 avss.n138 117.001
R327 avss.n163 avss.n155 117.001
R328 avss.n155 avss.n154 117.001
R329 avss.n175 avss.n70 117.001
R330 avss.n178 avss.n175 117.001
R331 avss.n176 avss.n72 117.001
R332 avss.n177 avss.n176 117.001
R333 avss.n169 avss.n168 117.001
R334 avss.n168 avss.n167 117.001
R335 avss.n253 avss.n252 117.001
R336 avss.n254 avss.n253 117.001
R337 avss.n116 avss.n115 117.001
R338 avss.n115 avss.n114 117.001
R339 avss.n103 avss.n96 117.001
R340 avss.n113 avss.n96 117.001
R341 avss.n100 avss.n45 117.001
R342 avss.n100 avss.n99 117.001
R343 avss.n52 avss.n47 117.001
R344 avss.n98 avss.n52 117.001
R345 avss.n56 avss.n53 117.001
R346 avss.n130 avss.n53 117.001
R347 avss.n59 avss.n57 117.001
R348 avss.n131 avss.n59 117.001
R349 avss.n64 avss.n60 117.001
R350 avss.n142 avss.n60 117.001
R351 avss.n157 avss.n144 117.001
R352 avss.n144 avss.n143 117.001
R353 avss.n147 avss.n145 117.001
R354 avss.n153 avss.n145 117.001
R355 avss.n150 avss.n148 117.001
R356 avss.n154 avss.n150 117.001
R357 avss.n151 avss.n69 117.001
R358 avss.n178 avss.n151 117.001
R359 avss.n75 avss.n71 117.001
R360 avss.n177 avss.n75 117.001
R361 avss.n79 avss.n76 117.001
R362 avss.n167 avss.n76 117.001
R363 avss.n82 avss.n80 117.001
R364 avss.n166 avss.n82 117.001
R365 avss.n83 avss.n81 117.001
R366 avss.n84 avss.n83 117.001
R367 avss.n267 avss.n266 117.001
R368 avss.n21 avss.n17 117.001
R369 avss.n21 avss.n11 117.001
R370 avss.n279 avss.n278 117.001
R371 avss.n280 avss.n279 117.001
R372 avss.n20 avss.n19 117.001
R373 avss.t44 avss.n263 114.418
R374 avss.n14 avss.t16 110.406
R375 avss.n99 avss.t138 101.523
R376 avss.n170 avss.n169 98.8418
R377 avss.t70 avss.n177 97.4624
R378 avss.t23 avss.n289 96.4472
R379 avss.t106 avss.n153 93.4015
R380 avss.n264 avss.t57 91.9439
R381 avss.t50 avss.t110 90.3558
R382 avss.n131 avss.t126 89.3406
R383 avss.t90 avss.t29 86.2949
R384 avss.n84 avss.t64 85.2797
R385 avss.t24 avss.n33 84.2645
R386 avss.t128 avss.n84 83.2492
R387 avss.n259 avss.n28 82.4476
R388 avss.t90 avss.t82 82.234
R389 avss.n252 avss.n36 82.0711
R390 avss.n111 avss.n40 82.0711
R391 avss.n219 avss.n80 82.0711
R392 avss.n85 avss.n80 82.0711
R393 avss.n162 avss.n148 82.0711
R394 avss.n163 avss.n162 82.0711
R395 avss.n226 avss.n69 82.0711
R396 avss.n226 avss.n70 82.0711
R397 avss.n158 avss.n157 82.0711
R398 avss.n158 avss.n135 82.0711
R399 avss.n161 avss.n147 82.0711
R400 avss.n161 avss.n156 82.0711
R401 avss.n63 avss.n57 82.0711
R402 avss.n133 avss.n63 82.0711
R403 avss.n65 avss.n64 82.0711
R404 avss.n134 avss.n65 82.0711
R405 avss.n242 avss.n47 82.0711
R406 avss.n242 avss.n48 82.0711
R407 avss.n127 avss.n56 82.0711
R408 avss.n128 avss.n127 82.0711
R409 avss.n103 avss.n102 82.0711
R410 avss.n102 avss.n101 82.0711
R411 avss.n243 avss.n45 82.0711
R412 avss.n243 avss.n46 82.0711
R413 avss.n116 avss.n40 82.0711
R414 avss.n220 avss.n79 82.0711
R415 avss.n165 avss.n79 82.0711
R416 avss.n78 avss.n71 82.0711
R417 avss.n225 avss.n71 82.0711
R418 avss.n225 avss.n72 82.0711
R419 avss.n169 avss.n165 82.0711
R420 avss.n108 avss.n36 81.6946
R421 avss.n111 avss.n110 81.6946
R422 avss.n182 avss.n148 81.6946
R423 avss.n164 avss.n163 81.6946
R424 avss.n149 avss.n69 81.6946
R425 avss.n172 avss.n70 81.6946
R426 avss.n157 avss.n146 81.6946
R427 avss.n188 avss.n135 81.6946
R428 avss.n183 avss.n147 81.6946
R429 avss.n156 avss.n136 81.6946
R430 avss.n236 avss.n57 81.6946
R431 avss.n191 avss.n133 81.6946
R432 avss.n64 avss.n58 81.6946
R433 avss.n189 avss.n134 81.6946
R434 avss.n55 avss.n47 81.6946
R435 avss.n125 avss.n48 81.6946
R436 avss.n237 avss.n56 81.6946
R437 avss.n192 avss.n128 81.6946
R438 avss.n118 avss.n103 81.6946
R439 avss.n101 avss.n91 81.6946
R440 avss.n119 avss.n45 81.6946
R441 avss.n124 avss.n46 81.6946
R442 avss.n117 avss.n116 81.6946
R443 avss.n171 avss.n72 81.6946
R444 avss.t83 avss.n254 81.2188
R445 avss.n107 avss.n28 80.9417
R446 avss.n131 avss.t124 79.1883
R447 avss.t50 avss.t112 78.1731
R448 avss.n264 avss.t121 77.6415
R449 avss.n282 avss.n281 75.7785
R450 avss.n153 avss.t55 75.1274
R451 avss.n288 avss.t123 75.0507
R452 avss.n265 avss.t51 72.4295
R453 avss.t102 avss.n274 72.4295
R454 avss.n289 avss.t2 72.0817
R455 avss.n177 avss.t105 71.0665
R456 avss.n108 avss.n107 70.0382
R457 avss.n99 avss.t118 67.0056
R458 avss.n265 avss.n15 66.7478
R459 avss.n274 avss.n273 66.7478
R460 avss.n199 avss.n198 65.9697
R461 avss.n263 avss.t75 55.1665
R462 avss.n276 avss.n19 50.3092
R463 avss.n267 avss.n18 50.106
R464 avss.n261 avss.n260 43.1857
R465 avss.t126 avss.n130 42.6401
R466 avss.n218 avss.n81 41.346
R467 avss.t48 avss.n256 40.8642
R468 avss.n268 avss.n267 40.4775
R469 avss.n106 avss.n105 39.9597
R470 avss.n23 avss.n19 39.8117
R471 avss.t96 avss.t31 39.5944
R472 avss.n154 avss.t106 38.5792
R473 avss.t46 avss.t7 35.5335
R474 avss.n178 avss.t70 34.5183
R475 avss.t94 avss.t37 31.4726
R476 avss.t138 avss.n98 30.4574
R477 avss.n113 avss.t9 28.4269
R478 avss.n214 avss.n81 27.9126
R479 avss.t88 avss.t10 27.4117
R480 avss.n105 avss.n27 25.3701
R481 avss.n261 avss.n27 25.361
R482 avss.n167 avss.t107 24.366
R483 avss.n277 avss.n276 23.6684
R484 avss.n277 avss.n18 23.4269
R485 avss.t33 avss.t113 23.3508
R486 avss.n143 avss.t134 20.3051
R487 avss.t6 avss.t86 19.2898
R488 avss.n258 avss.n27 17.4857
R489 avss.n117 avss.n38 17.1477
R490 avss.n120 avss.n118 17.1477
R491 avss.n120 avss.n119 17.1477
R492 avss.n238 avss.n55 17.1477
R493 avss.n238 avss.n237 17.1477
R494 avss.n236 avss.n235 17.1477
R495 avss.n235 avss.n58 17.1477
R496 avss.n184 avss.n146 17.1477
R497 avss.n184 avss.n183 17.1477
R498 avss.n182 avss.n181 17.1477
R499 avss.n181 avss.n149 17.1477
R500 avss.n107 avss.n106 17.1477
R501 avss.n109 avss.n108 17.1477
R502 avss.n110 avss.n109 17.1477
R503 avss.n123 avss.n91 17.1477
R504 avss.n124 avss.n123 17.1477
R505 avss.n126 avss.n125 17.1477
R506 avss.n191 avss.n190 17.1477
R507 avss.n190 avss.n189 17.1477
R508 avss.n188 avss.n187 17.1477
R509 avss.n187 avss.n136 17.1477
R510 avss.n173 avss.n164 17.1477
R511 avss.n173 avss.n172 17.1477
R512 avss.n171 avss.n170 17.1477
R513 avss.n219 avss.n218 17.0405
R514 avss.n221 avss.n78 17.0405
R515 avss.n221 avss.n220 17.0405
R516 avss.n215 avss.n85 16.8301
R517 avss.n225 avss.n224 16.8301
R518 avss.n287 avss.n286 16.7148
R519 avss.n12 avss.n8 16.7148
R520 avss.n291 avss.n290 16.7148
R521 avss.n201 avss.n200 16.7148
R522 avss.n162 avss.n68 16.6249
R523 avss.n159 avss.n158 16.6249
R524 avss.n232 avss.n63 16.6249
R525 avss.n242 avss.n241 16.6249
R526 avss.n102 avss.n44 16.6249
R527 avss.n142 avss.t133 16.2442
R528 avss.n251 avss.n38 15.7791
R529 avss.n278 avss.n277 15.7042
R530 avss.n260 avss.n259 15.6805
R531 avss.n251 avss.n250 15.2981
R532 avss.n259 avss.n258 15.2981
R533 avss.n272 avss.n271 15.1138
R534 avss.n271 avss.n269 14.9595
R535 avss.n193 avss.n126 14.6521
R536 avss.n270 avss.n17 13.6894
R537 avss.n202 avss.n201 13.3619
R538 avss.n215 avss.n214 12.7033
R539 avss.n166 avss.t84 12.1832
R540 avss.n292 avss.n291 11.4429
R541 avss.n118 avss.n117 10.4659
R542 avss.n119 avss.n55 10.4659
R543 avss.n237 avss.n236 10.4659
R544 avss.n146 avss.n58 10.4659
R545 avss.n183 avss.n182 10.4659
R546 avss.n110 avss.n91 10.4659
R547 avss.n125 avss.n124 10.4659
R548 avss.n192 avss.n191 10.4659
R549 avss.n189 avss.n188 10.4659
R550 avss.n164 avss.n136 10.4659
R551 avss.n172 avss.n171 10.4659
R552 avss.n149 avss.n78 10.4574
R553 avss.n220 avss.n219 10.4488
R554 avss.n224 avss.n74 10.4301
R555 avss.n165 avss.n85 10.4152
R556 avss.n226 avss.n225 10.3988
R557 avss.n162 avss.n161 10.3825
R558 avss.n158 avss.n65 10.3825
R559 avss.n127 avss.n63 10.3825
R560 avss.n243 avss.n242 10.3825
R561 avss.n102 avss.n40 10.3825
R562 avss.n227 avss.n68 10.3029
R563 avss.n160 avss.n159 10.3029
R564 avss.n232 avss.n231 10.3029
R565 avss.n241 avss.n51 10.3029
R566 avss.n244 avss.n44 10.3029
R567 avss.n250 avss.n249 10.3029
R568 avss.n37 avss.n29 9.81158
R569 avss.n195 avss.n194 9.70027
R570 avss.n208 avss.n194 9.38309
R571 avss.n211 avss.n90 8.52976
R572 avss.n114 avss.t68 8.12233
R573 avss.t87 avss.t127 7.15165
R574 avss.n165 avss.n74 6.4005
R575 avss.n227 avss.n226 6.32245
R576 avss.n161 avss.n160 6.32245
R577 avss.n231 avss.n65 6.32245
R578 avss.n127 avss.n51 6.32245
R579 avss.n244 avss.n243 6.32245
R580 avss.n249 avss.n40 6.32245
R581 avss.n252 avss.n37 4.88071
R582 avss.n7 avss.n5 4.00735
R583 avss.n13 avss.n5 4.00735
R584 avss.n285 avss.n6 4.00735
R585 avss.n13 avss.n6 4.00735
R586 avss.n4 avss.n2 4.00735
R587 avss.n33 avss.n4 4.00735
R588 avss.n198 avss.n3 4.00735
R589 avss.n33 avss.n3 4.00735
R590 avss.n271 avss.n270 3.79309
R591 avss.n254 avss.n33 3.04619
R592 avss.n193 avss.n192 2.4961
R593 avss.n41 avss.n37 2.3284
R594 avss.n214 avss.n213 2.3255
R595 avss.n23 avss.n22 2.3255
R596 avss.n268 avss.n10 2.3255
R597 avss.n89 avss 2.08383
R598 avss.n272 avss.n23 1.38845
R599 avss.n228 avss.n227 1.163
R600 avss.n160 avss.n66 1.163
R601 avss.n231 avss.n230 1.163
R602 avss.n51 avss.n50 1.163
R603 avss.n245 avss.n244 1.163
R604 avss.n249 avss.n248 1.163
R605 avss.n86 avss.n74 1.163
R606 avss.n213 avss.n212 1.1255
R607 avss.n270 avss.n9 1.03383
R608 avss.n269 avss.n268 0.925801
R609 avss.n293 avss.n292 0.885206
R610 avss.n203 avss.n202 0.885206
R611 avss.n207 avss.n1 0.577925
R612 avss.n199 avss.n197 0.577925
R613 avss.n42 avss.n41 0.570597
R614 avss.n87 avss.n86 0.563
R615 avss.n248 avss.n247 0.563
R616 avss.n246 avss.n245 0.563
R617 avss.n50 avss.n43 0.563
R618 avss.n230 avss.n229 0.563
R619 avss.n229 avss.n66 0.563
R620 avss.n229 avss.n228 0.563
R621 avss.n284 avss.n283 0.4655
R622 avss.n204 avss.n203 0.440907
R623 avss.n210 avss.n209 0.401201
R624 avss.n252 avss.n251 0.287571
R625 avss.n212 avss.n87 0.243877
R626 avss.n206 avss.n205 0.23753
R627 avss.n247 avss.n246 0.230632
R628 avss.n246 avss.n43 0.230632
R629 avss.n67 avss.n43 0.204142
R630 avss.n210 avss.n0 0.198
R631 avss.n205 avss.n196 0.184322
R632 avss.n194 avss.n193 0.173003
R633 avss.n259 avss.n29 0.163374
R634 avss.n195 avss.n42 0.146218
R635 avss.n211 avss.n210 0.128227
R636 avss.n278 avss.n17 0.119019
R637 avss.n204 avss.n197 0.115398
R638 avss.n206 avss.n0 0.107946
R639 avss.n205 avss.n204 0.10694
R640 avss.n247 avss.n42 0.104391
R641 avss.n197 avss.n196 0.0932734
R642 avss.n207 avss.n206 0.0927996
R643 avss.n90 avss.n89 0.068442
R644 avss.n293 avss.n0 0.0602048
R645 avss.n22 avss.n9 0.048994
R646 avss.n209 avss.n67 0.0428448
R647 avss avss.n293 0.0414213
R648 avss.n89 avss 0.0334815
R649 avss.n282 avss.n10 0.0319759
R650 avss.n87 avss.n67 0.0307152
R651 avss.n88 avss.n10 0.0164639
R652 avss.n283 avss.n9 0.0161626
R653 avss.n212 avss.n211 0.0108477
R654 avss.n208 avss.n207 0.0102951
R655 avss.n90 avss.n88 0.0068253
R656 avss.n209 avss.n208 0.0060003
R657 avss.n203 avss 0.00575492
R658 avss.n196 avss.n195 0.00372284
R659 avss.n229 avss.n67 0.00298644
R660 avss.n283 avss.n282 0.000650602
R661 a_1538_5653.n1 a_1538_5653.t3 660.701
R662 a_1538_5653.n0 a_1538_5653.t5 660.514
R663 a_1538_5653.n0 a_1538_5653.t7 660.466
R664 a_1538_5653.n0 a_1538_5653.t11 660.24
R665 a_1538_5653.n0 a_1538_5653.t12 660.24
R666 a_1538_5653.n1 a_1538_5653.t9 660.24
R667 a_1538_5653.t1 a_1538_5653.n1 660.24
R668 a_1538_5653.n0 a_1538_5653.t13 236.429
R669 a_1538_5653.n0 a_1538_5653.t4 212.572
R670 a_1538_5653.n0 a_1538_5653.t10 106.373
R671 a_1538_5653.n0 a_1538_5653.t17 106.373
R672 a_1538_5653.n0 a_1538_5653.t16 106.373
R673 a_1538_5653.n0 a_1538_5653.t18 106.373
R674 a_1538_5653.n0 a_1538_5653.t14 106.373
R675 a_1538_5653.n0 a_1538_5653.t15 106.373
R676 a_1538_5653.n0 a_1538_5653.t6 106.338
R677 a_1538_5653.n1 a_1538_5653.t0 106.338
R678 a_1538_5653.n1 a_1538_5653.t8 106.337
R679 a_1538_5653.n1 a_1538_5653.t2 106.335
R680 a_1538_5653.n1 a_1538_5653.n0 16.482
R681 avdd.n266 avdd.n23 28387.9
R682 avdd.n266 avdd.n265 28387.9
R683 avdd.n272 avdd.n23 19593
R684 avdd.n265 avdd.n264 19590.1
R685 avdd.n267 avdd.n26 15171.2
R686 avdd.n267 avdd.n24 15171.2
R687 avdd.n271 avdd.n24 10578.9
R688 avdd.n263 avdd.n26 10577.4
R689 avdd.n264 avdd.n22 6697.21
R690 avdd.n273 avdd.n272 6682.45
R691 avdd.n274 avdd.n22 5770.81
R692 avdd.n263 avdd.n20 3845.19
R693 avdd.n271 avdd.n21 3837.49
R694 avdd.n275 avdd.n21 3586.38
R695 avdd.n275 avdd.n20 3580.22
R696 avdd.n274 avdd.n273 3192.24
R697 avdd.n269 avdd.n268 1098.08
R698 avdd.n147 avdd.n130 1006.34
R699 avdd.n147 avdd.n131 1006.34
R700 avdd.n146 avdd.n130 1006.34
R701 avdd.n146 avdd.n131 1006.34
R702 avdd.n27 avdd.n25 881.597
R703 avdd.n210 avdd.n73 841.241
R704 avdd.n210 avdd.n74 841.241
R705 avdd.n74 avdd.n72 841.241
R706 avdd.n73 avdd.n72 841.241
R707 avdd.n203 avdd.n78 841.241
R708 avdd.n203 avdd.n79 841.241
R709 avdd.n202 avdd.n79 841.241
R710 avdd.n202 avdd.n78 841.241
R711 avdd.n187 avdd.n95 841.241
R712 avdd.n187 avdd.n96 841.241
R713 avdd.n96 avdd.n94 841.241
R714 avdd.n95 avdd.n94 841.241
R715 avdd.n173 avdd.n109 841.241
R716 avdd.n173 avdd.n110 841.241
R717 avdd.n110 avdd.n103 841.241
R718 avdd.n109 avdd.n103 841.241
R719 avdd.n152 avdd.n125 841.241
R720 avdd.n153 avdd.n125 841.241
R721 avdd.n166 avdd.n115 841.241
R722 avdd.n165 avdd.n115 841.241
R723 avdd.n70 avdd.n68 841.241
R724 avdd.n211 avdd.n68 841.241
R725 avdd.n211 avdd.n67 841.241
R726 avdd.n70 avdd.n67 841.241
R727 avdd.n194 avdd.n81 841.241
R728 avdd.n194 avdd.n82 841.241
R729 avdd.n85 avdd.n82 841.241
R730 avdd.n85 avdd.n81 841.241
R731 avdd.n92 avdd.n90 841.241
R732 avdd.n188 avdd.n90 841.241
R733 avdd.n188 avdd.n89 841.241
R734 avdd.n92 avdd.n89 841.241
R735 avdd.n174 avdd.n105 841.241
R736 avdd.n107 avdd.n105 841.241
R737 avdd.n107 avdd.n104 841.241
R738 avdd.n174 avdd.n104 841.241
R739 avdd.n122 avdd.n117 841.241
R740 avdd.n122 avdd.n118 841.241
R741 avdd.n135 avdd.n118 841.241
R742 avdd.n135 avdd.n117 841.241
R743 avdd.n246 avdd.n42 841.241
R744 avdd.n247 avdd.n42 841.241
R745 avdd.n230 avdd.n225 841.241
R746 avdd.n225 avdd.n224 841.241
R747 avdd.n45 avdd.n40 841.241
R748 avdd.n222 avdd.n220 841.241
R749 avdd.n231 avdd.n220 841.241
R750 avdd.n46 avdd.n45 841.241
R751 avdd.n301 avdd.n6 841.241
R752 avdd.n301 avdd.n7 841.241
R753 avdd.n297 avdd.n7 841.241
R754 avdd.n297 avdd.n6 841.241
R755 avdd.n295 avdd.n11 841.241
R756 avdd.n295 avdd.n12 841.241
R757 avdd.n286 avdd.n12 841.241
R758 avdd.n286 avdd.n11 841.241
R759 avdd.n305 avdd.n4 841.241
R760 avdd.n306 avdd.n4 841.241
R761 avdd.n306 avdd.n3 841.241
R762 avdd.n305 avdd.n3 841.241
R763 avdd.n292 avdd.n13 841.241
R764 avdd.n292 avdd.n288 841.241
R765 avdd.n288 avdd.n14 841.241
R766 avdd.n14 avdd.n13 841.241
R767 avdd.n270 avdd.n269 823.929
R768 avdd.n159 avdd.t10 661.426
R769 avdd.n251 avdd.t28 660.576
R770 avdd.n251 avdd.t15 660.562
R771 avdd.n99 avdd.t2 660.562
R772 avdd.n36 avdd.t4 660.562
R773 avdd.n35 avdd.t6 660.562
R774 avdd.n158 avdd.t13 660.562
R775 avdd.n161 avdd.t16 660.562
R776 avdd.n289 avdd.t25 660.391
R777 avdd.n0 avdd.t29 660.38
R778 avdd.n237 avdd.t8 660.341
R779 avdd.n236 avdd.t11 660.34
R780 avdd.n237 avdd.t18 660.327
R781 avdd.n236 avdd.t19 660.319
R782 avdd.n262 avdd.n27 654.298
R783 avdd.n58 avdd.n53 422.587
R784 avdd.n58 avdd.n57 422.587
R785 avdd.n50 avdd.n48 422.587
R786 avdd.n50 avdd.n43 422.587
R787 avdd.n155 avdd.n114 422.587
R788 avdd.n155 avdd.n120 422.587
R789 avdd.n233 avdd.n219 422.587
R790 avdd.n233 avdd.n232 422.587
R791 avdd.n63 avdd.n61 422.587
R792 avdd.n63 avdd.n62 422.587
R793 avdd.n152 avdd.n114 418.656
R794 avdd.n166 avdd.n114 418.656
R795 avdd.n153 avdd.n120 418.656
R796 avdd.n165 avdd.n120 418.656
R797 avdd.n246 avdd.n48 418.656
R798 avdd.n242 avdd.n48 418.656
R799 avdd.n242 avdd.n53 418.656
R800 avdd.n230 avdd.n53 418.656
R801 avdd.n247 avdd.n43 418.656
R802 avdd.n241 avdd.n43 418.656
R803 avdd.n241 avdd.n57 418.656
R804 avdd.n224 avdd.n57 418.656
R805 avdd.n61 avdd.n40 418.656
R806 avdd.n61 avdd.n54 418.656
R807 avdd.n219 avdd.n54 418.656
R808 avdd.n222 avdd.n219 418.656
R809 avdd.n62 avdd.n46 418.656
R810 avdd.n62 avdd.n55 418.656
R811 avdd.n232 avdd.n55 418.656
R812 avdd.n232 avdd.n231 418.656
R813 avdd.n270 avdd.n18 282.248
R814 avdd.n261 avdd.n28 242.221
R815 avdd.n277 avdd.n276 175.579
R816 avdd.n133 avdd.n130 175.579
R817 avdd.n29 avdd.n19 171.523
R818 avdd.n274 avdd.n16 168.218
R819 avdd.t9 avdd.n126 149.226
R820 avdd.t9 avdd.n116 149.226
R821 avdd.t12 avdd.n116 149.226
R822 avdd.t12 avdd.n119 149.226
R823 avdd.t0 avdd.n106 149.226
R824 avdd.t0 avdd.n108 149.226
R825 avdd.t1 avdd.n91 149.226
R826 avdd.t1 avdd.n93 149.226
R827 avdd.t3 avdd.n80 149.226
R828 avdd.t3 avdd.n83 149.226
R829 avdd.t5 avdd.n69 149.226
R830 avdd.t5 avdd.n71 149.226
R831 avdd.t14 avdd.n44 149.226
R832 avdd.t14 avdd.n47 149.226
R833 avdd.t7 avdd.n47 149.226
R834 avdd.t7 avdd.n56 149.226
R835 avdd.t17 avdd.n56 149.226
R836 avdd.t17 avdd.n223 149.226
R837 avdd.n133 avdd.n132 149.161
R838 avdd.n119 avdd.n106 133.113
R839 avdd.n108 avdd.n91 133.113
R840 avdd.n93 avdd.n80 133.113
R841 avdd.n83 avdd.n69 133.113
R842 avdd.n71 avdd.n44 133.113
R843 avdd.t23 avdd.n5 128.886
R844 avdd.t23 avdd.n8 128.886
R845 avdd.t24 avdd.n287 125.255
R846 avdd.n293 avdd.t26 125.255
R847 avdd.n294 avdd.n5 111.338
R848 avdd.n144 avdd.n134 106.541
R849 avdd.n198 avdd.n197 91.9447
R850 avdd.n86 avdd.n84 91.9447
R851 avdd.n179 avdd.n178 91.9447
R852 avdd.n136 avdd.n121 91.9447
R853 avdd.n249 avdd.n39 91.9447
R854 avdd.n139 avdd.n102 91.9447
R855 avdd.n132 avdd.n126 91.0772
R856 avdd.n162 avdd.n111 90.0623
R857 avdd.n199 avdd.n75 90.0623
R858 avdd.n182 avdd.n181 90.0623
R859 avdd.n177 avdd.n98 90.0623
R860 avdd.n157 avdd.n156 90.0623
R861 avdd.n250 avdd.n38 90.0623
R862 avdd.n65 avdd.n37 85.4593
R863 avdd.n200 avdd.n195 85.4593
R864 avdd.n183 avdd.n87 85.4593
R865 avdd.n176 avdd.n101 85.4593
R866 avdd.n163 avdd.n123 85.4593
R867 avdd.n235 avdd.n234 85.4593
R868 avdd.n64 avdd.n41 85.4593
R869 avdd.n213 avdd.n65 85.0829
R870 avdd.n197 avdd.n66 85.0829
R871 avdd.n195 avdd.n193 85.0829
R872 avdd.n191 avdd.n86 85.0829
R873 avdd.n190 avdd.n87 85.0829
R874 avdd.n178 avdd.n88 85.0829
R875 avdd.n137 avdd.n101 85.0829
R876 avdd.n143 avdd.n136 85.0829
R877 avdd.n141 avdd.n123 85.0829
R878 avdd.n234 avdd.n218 85.0829
R879 avdd.n214 avdd.n39 85.0829
R880 avdd.n216 avdd.n64 85.0829
R881 avdd.n140 avdd.n139 85.0829
R882 avdd.n51 avdd.n41 83.9534
R883 avdd.n207 avdd.n37 83.9534
R884 avdd.n200 avdd.n76 83.9534
R885 avdd.n184 avdd.n183 83.9534
R886 avdd.n176 avdd.n100 83.9534
R887 avdd.n163 avdd.n112 83.9534
R888 avdd.n127 avdd.n124 83.9534
R889 avdd.n235 avdd.n59 83.577
R890 avdd.n59 avdd.n52 82.824
R891 avdd.n244 avdd.n51 82.824
R892 avdd.n169 avdd.n111 82.824
R893 avdd.n208 avdd.n207 82.824
R894 avdd.n206 avdd.n75 82.824
R895 avdd.n205 avdd.n76 82.824
R896 avdd.n181 avdd.n77 82.824
R897 avdd.n185 avdd.n184 82.824
R898 avdd.n170 avdd.n98 82.824
R899 avdd.n171 avdd.n100 82.824
R900 avdd.n156 avdd.n113 82.824
R901 avdd.n168 avdd.n112 82.824
R902 avdd.n150 avdd.n127 82.824
R903 avdd.n49 avdd.n38 82.824
R904 avdd.n134 avdd.n129 64.7534
R905 avdd.n149 avdd.n128 57.1448
R906 avdd.n229 avdd.n228 54.5383
R907 avdd.n285 avdd.n10 51.1301
R908 avdd.n302 avdd.n300 50.4217
R909 avdd.n268 avdd.n25 49.7553
R910 avdd.n145 avdd.n128 49.2624
R911 avdd.n164 avdd.n117 46.2505
R912 avdd.t12 avdd.n117 46.2505
R913 avdd.n175 avdd.n174 46.2505
R914 avdd.n174 avdd.t0 46.2505
R915 avdd.n180 avdd.n92 46.2505
R916 avdd.t1 avdd.n92 46.2505
R917 avdd.n201 avdd.n81 46.2505
R918 avdd.t3 avdd.n81 46.2505
R919 avdd.n196 avdd.n70 46.2505
R920 avdd.t5 avdd.n70 46.2505
R921 avdd.n165 avdd.n164 46.2505
R922 avdd.t12 avdd.n165 46.2505
R923 avdd.n175 avdd.n103 46.2505
R924 avdd.t0 avdd.n103 46.2505
R925 avdd.n180 avdd.n94 46.2505
R926 avdd.t1 avdd.n94 46.2505
R927 avdd.n202 avdd.n201 46.2505
R928 avdd.t3 avdd.n202 46.2505
R929 avdd.n196 avdd.n72 46.2505
R930 avdd.t5 avdd.n72 46.2505
R931 avdd.n148 avdd.n147 46.2505
R932 avdd.n147 avdd.t27 46.2505
R933 avdd.n154 avdd.n153 46.2505
R934 avdd.n153 avdd.t9 46.2505
R935 avdd.n167 avdd.n166 46.2505
R936 avdd.n166 avdd.t12 46.2505
R937 avdd.n152 avdd.n151 46.2505
R938 avdd.t9 avdd.n152 46.2505
R939 avdd.n173 avdd.n172 46.2505
R940 avdd.t0 avdd.n173 46.2505
R941 avdd.n187 avdd.n186 46.2505
R942 avdd.t1 avdd.n187 46.2505
R943 avdd.n204 avdd.n203 46.2505
R944 avdd.n203 avdd.t3 46.2505
R945 avdd.n210 avdd.n209 46.2505
R946 avdd.t5 avdd.n210 46.2505
R947 avdd.n230 avdd.n229 46.2505
R948 avdd.t17 avdd.n230 46.2505
R949 avdd.n243 avdd.n242 46.2505
R950 avdd.n242 avdd.t7 46.2505
R951 avdd.n246 avdd.n245 46.2505
R952 avdd.t14 avdd.n246 46.2505
R953 avdd.n241 avdd.n240 46.2505
R954 avdd.t7 avdd.n241 46.2505
R955 avdd.n224 avdd.n60 46.2505
R956 avdd.t17 avdd.n224 46.2505
R957 avdd.n222 avdd.n60 46.2505
R958 avdd.t17 avdd.n222 46.2505
R959 avdd.n240 avdd.n54 46.2505
R960 avdd.t7 avdd.n54 46.2505
R961 avdd.n231 avdd.n221 46.2505
R962 avdd.n231 avdd.t17 46.2505
R963 avdd.n217 avdd.n55 46.2505
R964 avdd.t7 avdd.n55 46.2505
R965 avdd.n248 avdd.n40 46.2505
R966 avdd.t14 avdd.n40 46.2505
R967 avdd.n248 avdd.n247 46.2505
R968 avdd.n247 avdd.t14 46.2505
R969 avdd.n142 avdd.n118 46.2505
R970 avdd.t12 avdd.n118 46.2505
R971 avdd.n138 avdd.n107 46.2505
R972 avdd.t0 avdd.n107 46.2505
R973 avdd.n189 avdd.n188 46.2505
R974 avdd.n188 avdd.t1 46.2505
R975 avdd.n192 avdd.n82 46.2505
R976 avdd.t3 avdd.n82 46.2505
R977 avdd.n212 avdd.n211 46.2505
R978 avdd.n211 avdd.t5 46.2505
R979 avdd.n215 avdd.n46 46.2505
R980 avdd.t14 avdd.n46 46.2505
R981 avdd.n146 avdd.n145 46.2505
R982 avdd.t27 avdd.n146 46.2505
R983 avdd.n283 avdd.n13 46.2505
R984 avdd.t24 avdd.n13 46.2505
R985 avdd.n288 avdd.n15 46.2505
R986 avdd.n288 avdd.t24 46.2505
R987 avdd.n305 avdd.n304 46.2505
R988 avdd.t23 avdd.n305 46.2505
R989 avdd.n307 avdd.n306 46.2505
R990 avdd.n306 avdd.t23 46.2505
R991 avdd.n11 avdd.n10 46.2505
R992 avdd.t26 avdd.n11 46.2505
R993 avdd.n282 avdd.n12 46.2505
R994 avdd.t26 avdd.n12 46.2505
R995 avdd.n300 avdd.n6 46.2505
R996 avdd.t23 avdd.n6 46.2505
R997 avdd.n304 avdd.n7 46.2505
R998 avdd.t23 avdd.n7 46.2505
R999 avdd.n144 avdd.n143 44.7603
R1000 avdd.n255 avdd.t21 43.8338
R1001 avdd.n32 avdd.t22 42.394
R1002 avdd.n32 avdd.t20 42.3922
R1003 avdd.n277 avdd.n18 42.2199
R1004 avdd.n226 avdd.n221 40.8829
R1005 avdd.n150 avdd.n149 39.5172
R1006 avdd.n136 avdd.n135 37.0005
R1007 avdd.n135 avdd.n116 37.0005
R1008 avdd.n123 avdd.n122 37.0005
R1009 avdd.n122 avdd.n119 37.0005
R1010 avdd.n105 avdd.n101 37.0005
R1011 avdd.n108 avdd.n105 37.0005
R1012 avdd.n178 avdd.n89 37.0005
R1013 avdd.n91 avdd.n89 37.0005
R1014 avdd.n90 avdd.n87 37.0005
R1015 avdd.n93 avdd.n90 37.0005
R1016 avdd.n86 avdd.n85 37.0005
R1017 avdd.n85 avdd.n80 37.0005
R1018 avdd.n195 avdd.n194 37.0005
R1019 avdd.n194 avdd.n83 37.0005
R1020 avdd.n197 avdd.n67 37.0005
R1021 avdd.n69 avdd.n67 37.0005
R1022 avdd.n68 avdd.n65 37.0005
R1023 avdd.n71 avdd.n68 37.0005
R1024 avdd.n156 avdd.n155 37.0005
R1025 avdd.n155 avdd.n116 37.0005
R1026 avdd.n115 avdd.n112 37.0005
R1027 avdd.n119 avdd.n115 37.0005
R1028 avdd.n111 avdd.n109 37.0005
R1029 avdd.n109 avdd.n106 37.0005
R1030 avdd.n110 avdd.n100 37.0005
R1031 avdd.n110 avdd.n108 37.0005
R1032 avdd.n98 avdd.n95 37.0005
R1033 avdd.n95 avdd.n91 37.0005
R1034 avdd.n184 avdd.n96 37.0005
R1035 avdd.n96 avdd.n93 37.0005
R1036 avdd.n181 avdd.n78 37.0005
R1037 avdd.n80 avdd.n78 37.0005
R1038 avdd.n79 avdd.n76 37.0005
R1039 avdd.n83 avdd.n79 37.0005
R1040 avdd.n75 avdd.n73 37.0005
R1041 avdd.n73 avdd.n69 37.0005
R1042 avdd.n207 avdd.n74 37.0005
R1043 avdd.n74 avdd.n71 37.0005
R1044 avdd.n51 avdd.n50 37.0005
R1045 avdd.n50 avdd.n47 37.0005
R1046 avdd.n59 avdd.n58 37.0005
R1047 avdd.n58 avdd.n56 37.0005
R1048 avdd.n127 avdd.n125 37.0005
R1049 avdd.n126 avdd.n125 37.0005
R1050 avdd.n42 avdd.n38 37.0005
R1051 avdd.n44 avdd.n42 37.0005
R1052 avdd.n228 avdd.n225 37.0005
R1053 avdd.n225 avdd.n223 37.0005
R1054 avdd.n234 avdd.n233 37.0005
R1055 avdd.n233 avdd.n56 37.0005
R1056 avdd.n226 avdd.n220 37.0005
R1057 avdd.n223 avdd.n220 37.0005
R1058 avdd.n45 avdd.n39 37.0005
R1059 avdd.n45 avdd.n44 37.0005
R1060 avdd.n64 avdd.n63 37.0005
R1061 avdd.n63 avdd.n47 37.0005
R1062 avdd.n139 avdd.n104 37.0005
R1063 avdd.n106 avdd.n104 37.0005
R1064 avdd.n281 avdd.n14 37.0005
R1065 avdd.n16 avdd.n14 37.0005
R1066 avdd.n292 avdd.n291 37.0005
R1067 avdd.n293 avdd.n292 37.0005
R1068 avdd.n291 avdd.n3 37.0005
R1069 avdd.n5 avdd.n3 37.0005
R1070 avdd.n4 avdd.n1 37.0005
R1071 avdd.n8 avdd.n4 37.0005
R1072 avdd.n286 avdd.n285 37.0005
R1073 avdd.n287 avdd.n286 37.0005
R1074 avdd.n296 avdd.n295 37.0005
R1075 avdd.n295 avdd.n294 37.0005
R1076 avdd.n298 avdd.n297 37.0005
R1077 avdd.n297 avdd.n5 37.0005
R1078 avdd.n302 avdd.n301 37.0005
R1079 avdd.n301 avdd.n8 37.0005
R1080 avdd.n243 avdd.n52 36.3525
R1081 avdd.n229 avdd.n52 36.3525
R1082 avdd.n275 avdd.n274 35.604
R1083 avdd.n130 avdd.n128 31.0027
R1084 avdd.n148 avdd.n129 29.6145
R1085 avdd.n308 avdd.n307 26.6196
R1086 avdd.n134 avdd.n131 26.4291
R1087 avdd.n132 avdd.n131 26.4291
R1088 avdd.n280 avdd.n15 25.9151
R1089 avdd.n29 avdd.n28 23.6252
R1090 avdd.n300 avdd.n299 23.2301
R1091 avdd.n299 avdd.n10 23.2301
R1092 avdd.n284 avdd.n281 23.1206
R1093 avdd.n303 avdd.n1 23.0608
R1094 avdd.n303 avdd.n302 23.0608
R1095 avdd.n281 avdd.n280 23.0608
R1096 avdd.n244 avdd.n243 22.7618
R1097 avdd.n285 avdd.n284 22.7005
R1098 avdd.n308 avdd.n1 21.9434
R1099 avdd.n307 avdd.n2 20.2328
R1100 avdd.n15 avdd.n2 20.2328
R1101 avdd.n291 avdd.n9 19.0862
R1102 avdd.n227 avdd.n226 18.6261
R1103 avdd.n228 avdd.n227 18.2979
R1104 avdd.n218 avdd.n217 17.3661
R1105 avdd.n221 avdd.n218 17.3661
R1106 avdd.n217 avdd.n216 17.2595
R1107 avdd.n151 avdd.n150 17.1477
R1108 avdd.n151 avdd.n113 17.1477
R1109 avdd.n167 avdd.n113 17.1477
R1110 avdd.n168 avdd.n167 17.1477
R1111 avdd.n172 avdd.n169 17.1477
R1112 avdd.n172 avdd.n171 17.1477
R1113 avdd.n186 avdd.n185 17.1477
R1114 avdd.n204 avdd.n77 17.1477
R1115 avdd.n205 avdd.n204 17.1477
R1116 avdd.n209 avdd.n206 17.1477
R1117 avdd.n209 avdd.n208 17.1477
R1118 avdd.n245 avdd.n49 17.1477
R1119 avdd.n245 avdd.n244 17.1477
R1120 avdd.n145 avdd.n144 17.1477
R1121 avdd.n143 avdd.n142 17.1477
R1122 avdd.n142 avdd.n141 17.1477
R1123 avdd.n140 avdd.n138 17.1477
R1124 avdd.n138 avdd.n137 17.1477
R1125 avdd.n189 avdd.n88 17.1477
R1126 avdd.n190 avdd.n189 17.1477
R1127 avdd.n192 avdd.n191 17.1477
R1128 avdd.n193 avdd.n192 17.1477
R1129 avdd.n212 avdd.n66 17.1477
R1130 avdd.n213 avdd.n212 17.1477
R1131 avdd.n215 avdd.n214 17.1477
R1132 avdd.n216 avdd.n215 17.1477
R1133 avdd.n299 avdd.n298 16.2647
R1134 avdd.n227 avdd.n60 15.383
R1135 avdd.n169 avdd.n168 15.2961
R1136 avdd.n171 avdd.n170 15.2961
R1137 avdd.n185 avdd.n77 15.2961
R1138 avdd.n206 avdd.n205 15.2961
R1139 avdd.n208 avdd.n49 15.2961
R1140 avdd.n141 avdd.n140 15.2961
R1141 avdd.n137 avdd.n88 15.2961
R1142 avdd.n191 avdd.n190 15.2961
R1143 avdd.n193 avdd.n66 15.2961
R1144 avdd.n214 avdd.n213 15.2961
R1145 avdd.n284 avdd.n283 15.193
R1146 avdd.n304 avdd.n303 14.8746
R1147 avdd.n296 avdd.n9 13.2702
R1148 avdd.n154 avdd.n124 12.0642
R1149 avdd.n196 avdd.n37 11.9584
R1150 avdd.n201 avdd.n200 11.9584
R1151 avdd.n183 avdd.n180 11.9584
R1152 avdd.n176 avdd.n175 11.9584
R1153 avdd.n164 avdd.n163 11.9584
R1154 avdd.n248 avdd.n41 11.9584
R1155 avdd.n235 avdd.n60 11.9542
R1156 avdd.n240 avdd.n41 11.9327
R1157 avdd.n304 avdd.n9 11.6153
R1158 avdd.n282 avdd.n9 11.365
R1159 avdd.n157 avdd.n154 11.0892
R1160 avdd.n186 avdd.n97 10.9489
R1161 avdd.n262 avdd.n261 10.3151
R1162 avdd.n239 avdd.n235 10.1175
R1163 avdd.n250 avdd.n37 9.77806
R1164 avdd.n200 avdd.n199 9.77806
R1165 avdd.n183 avdd.n182 9.77806
R1166 avdd.n177 avdd.n176 9.77806
R1167 avdd.n163 avdd.n162 9.77806
R1168 avdd.n291 avdd.n290 8.8005
R1169 avdd.n290 avdd.n2 7.6005
R1170 avdd.n129 avdd.n124 7.36333
R1171 avdd.n149 avdd.n148 7.12777
R1172 avdd.n28 avdd.n20 7.11588
R1173 avdd.n22 avdd.n20 7.11588
R1174 avdd.n21 avdd.n18 7.11588
R1175 avdd.n273 avdd.n21 7.11588
R1176 avdd.n170 avdd.n97 6.19924
R1177 avdd.n276 avdd.n275 4.74409
R1178 avdd.n263 avdd.n262 4.11161
R1179 avdd.n264 avdd.n263 4.11161
R1180 avdd.n271 avdd.n270 4.11161
R1181 avdd.n272 avdd.n271 4.11161
R1182 avdd.n287 avdd.n16 3.63107
R1183 avdd.t24 avdd.t26 3.63107
R1184 avdd.n294 avdd.n293 3.63107
R1185 avdd.n309 avdd.n308 3.10844
R1186 avdd.n280 avdd.n279 3.1005
R1187 avdd.n276 avdd.n19 2.57768
R1188 avdd.n240 avdd.n239 1.78915
R1189 avdd.n278 avdd.n277 1.43458
R1190 avdd.n268 avdd.n267 1.39148
R1191 avdd.n267 avdd.n266 1.39148
R1192 avdd.n30 avdd.n17 1.29749
R1193 avdd.n27 avdd.n26 1.1864
R1194 avdd.n265 avdd.n26 1.1864
R1195 avdd.n269 avdd.n24 1.1864
R1196 avdd.n24 avdd.n23 1.1864
R1197 avdd.n257 avdd.n32 1.03788
R1198 avdd.n290 avdd.n289 0.9305
R1199 avdd.n261 avdd.n260 0.885206
R1200 avdd.n256 avdd.n255 0.87315
R1201 avdd.n278 avdd.n17 0.863903
R1202 avdd.n199 avdd.n35 0.7755
R1203 avdd.n182 avdd.n36 0.7755
R1204 avdd.n177 avdd.n99 0.7755
R1205 avdd.n158 avdd.n157 0.7755
R1206 avdd.n239 avdd.n238 0.7755
R1207 avdd.n251 avdd.n250 0.7755
R1208 avdd.n162 avdd.n161 0.7755
R1209 avdd.n259 avdd.n30 0.640881
R1210 avdd.n30 avdd.n29 0.586059
R1211 avdd.n33 avdd.n31 0.553476
R1212 avdd.n259 avdd.n258 0.482723
R1213 avdd.n159 avdd.n158 0.376423
R1214 avdd.n161 avdd.n160 0.3755
R1215 avdd.n99 avdd.n34 0.3755
R1216 avdd.n252 avdd.n36 0.3755
R1217 avdd.n252 avdd.n35 0.3755
R1218 avdd.n252 avdd.n251 0.3755
R1219 avdd.n283 avdd.n282 0.359379
R1220 avdd.n198 avdd.n196 0.281202
R1221 avdd.n201 avdd.n84 0.281202
R1222 avdd.n180 avdd.n179 0.281202
R1223 avdd.n175 avdd.n102 0.281202
R1224 avdd.n164 avdd.n121 0.281202
R1225 avdd.n249 avdd.n248 0.281202
R1226 avdd.n255 avdd.n25 0.2618
R1227 avdd.n238 avdd.n237 0.250671
R1228 avdd.n257 avdd.n256 0.249606
R1229 avdd.n238 avdd.n236 0.249014
R1230 avdd.n160 avdd.n34 0.244171
R1231 avdd.n19 avdd.n17 0.233
R1232 avdd.n254 avdd.n33 0.220143
R1233 avdd.n97 avdd.n33 0.213887
R1234 avdd.n258 avdd.n31 0.206498
R1235 avdd.n258 avdd.n257 0.17749
R1236 avdd.n159 avdd.n31 0.165091
R1237 avdd.n253 avdd.n34 0.14963
R1238 avdd.n279 avdd.n0 0.122295
R1239 avdd.n160 avdd.n159 0.121149
R1240 avdd.n309 avdd.n0 0.119303
R1241 avdd.n298 avdd.n296 0.117931
R1242 avdd.n257 avdd.n254 0.113588
R1243 avdd.n260 avdd.n259 0.082678
R1244 avdd.n199 avdd.n198 0.0573889
R1245 avdd.n182 avdd.n84 0.0573889
R1246 avdd.n179 avdd.n177 0.0573889
R1247 avdd.n157 avdd.n121 0.0573889
R1248 avdd.n250 avdd.n249 0.0573889
R1249 avdd.n162 avdd.n102 0.0573889
R1250 avdd.n254 avdd.n253 0.0547069
R1251 avdd.t27 avdd.n133 0.0359565
R1252 avdd.n256 avdd 0.0256565
R1253 avdd.n279 avdd.n278 0.0139615
R1254 avdd avdd.n309 0.0139615
R1255 avdd.n260 avdd 0.0054195
R1256 avdd.n289 avdd.n0 0.00377715
R1257 avdd.n253 avdd.n252 0.000801568
R1258 ena.n4 ena.t1 396.2
R1259 ena.n4 ena.t2 381.825
R1260 ena.n0 ena.t5 305.348
R1261 ena.n2 ena.t4 196.596
R1262 ena.n1 ena.t3 112.246
R1263 ena.n1 ena.t0 110.207
R1264 ena.n4 ena.n3 4.5005
R1265 ena.n3 ena.n2 2.03668
R1266 ena.n3 ena.n0 1.72267
R1267 ena.n2 ena.n1 1.20571
R1268 ena.n0 ena 0.83638
R1269 ena ena.n4 0.062375
R1270 rc_osc_level_shifter_0.outb_h.n0 rc_osc_level_shifter_0.outb_h.t0 660.24
R1271 rc_osc_level_shifter_0.outb_h.n0 rc_osc_level_shifter_0.outb_h.t1 235.004
R1272 rc_osc_level_shifter_0.outb_h rc_osc_level_shifter_0.outb_h.t2 124.719
R1273 rc_osc_level_shifter_0.outb_h.n0 rc_osc_level_shifter_0.outb_h.t3 116.334
R1274 rc_osc_level_shifter_0.outb_h.n0 rc_osc_level_shifter_0.outb_h.t4 107.222
R1275 rc_osc_level_shifter_0.outb_h rc_osc_level_shifter_0.outb_h.n0 11.5134
R1276 dvdd.n25 dvdd.n24 1962.21
R1277 dvdd.n22 dvdd.n16 1796.47
R1278 dvdd.n16 dvdd.n15 1796.47
R1279 dvdd.n15 dvdd.n9 1796.47
R1280 dvdd.n36 dvdd.n5 1312.94
R1281 dvdd.n30 dvdd.n7 704.168
R1282 dvdd.n36 dvdd.n4 697.11
R1283 dvdd.n22 dvdd.n11 681.178
R1284 dvdd.n11 dvdd.n10 678.173
R1285 dvdd.n0 dvdd.t5 662.327
R1286 dvdd.n34 dvdd.n4 596.572
R1287 dvdd.n34 dvdd.n7 589.715
R1288 dvdd.n28 dvdd.n27 497.647
R1289 dvdd.n28 dvdd.n7 497.647
R1290 dvdd.n10 dvdd.n4 497.647
R1291 dvdd.n35 dvdd.t4 334.182
R1292 dvdd.n25 dvdd.t4 332.08
R1293 dvdd.t6 dvdd.n35 332.08
R1294 dvdd.n16 dvdd.t2 301.038
R1295 dvdd.n6 dvdd.n5 276.377
R1296 dvdd.n1 dvdd.t7 228.498
R1297 dvdd.n39 dvdd.t3 227.81
R1298 dvdd.n27 dvdd.n26 220.851
R1299 dvdd.n33 dvdd.n2 212.987
R1300 dvdd.n20 dvdd.n2 187.03
R1301 dvdd.n21 dvdd.n19 172.083
R1302 dvdd.n19 dvdd.n18 171.689
R1303 dvdd.n12 dvdd.t1 170.321
R1304 dvdd.n24 dvdd.t0 148.036
R1305 dvdd.n26 dvdd.n11 141.702
R1306 dvdd.n36 dvdd.t6 101.505
R1307 dvdd.n18 dvdd.n17 98.9414
R1308 dvdd.n10 dvdd.n2 92.5858
R1309 dvdd.n29 dvdd.n28 92.5005
R1310 dvdd.n28 dvdd.t4 92.5005
R1311 dvdd.n19 dvdd.n16 92.5005
R1312 dvdd.n17 dvdd.n9 92.5005
R1313 dvdd.n24 dvdd.n9 92.5005
R1314 dvdd.n31 dvdd.n30 92.5005
R1315 dvdd.n10 dvdd.t4 92.5005
R1316 dvdd.n37 dvdd.n36 92.5005
R1317 dvdd.n31 dvdd.n3 90.9905
R1318 dvdd.n30 dvdd.n6 77.441
R1319 dvdd.n32 dvdd.n31 75.1118
R1320 dvdd.n27 dvdd.n9 74.6438
R1321 dvdd.n33 dvdd.n32 62.9034
R1322 dvdd.n23 dvdd.t2 61.7891
R1323 dvdd.t0 dvdd.n23 61.7891
R1324 dvdd.n26 dvdd.n14 61.6672
R1325 dvdd.n26 dvdd.n25 61.6672
R1326 dvdd.n22 dvdd.n21 53.2393
R1327 dvdd.n32 dvdd.n29 53.0829
R1328 dvdd.n37 dvdd.n3 52.7584
R1329 dvdd.n29 dvdd.n8 50.824
R1330 dvdd.n23 dvdd.n22 46.2505
R1331 dvdd.n18 dvdd.n15 46.2505
R1332 dvdd.n23 dvdd.n15 46.2505
R1333 dvdd.n5 dvdd.n3 46.2505
R1334 dvdd.n34 dvdd.n33 46.2505
R1335 dvdd.n35 dvdd.n34 46.2505
R1336 dvdd.n21 dvdd.n20 31.463
R1337 dvdd.n38 dvdd.n2 27.0618
R1338 dvdd.t6 dvdd.n6 22.3157
R1339 dvdd.n14 dvdd.n13 18.5605
R1340 dvdd.n20 dvdd.n14 15.7445
R1341 dvdd.n17 dvdd.n8 4.0965
R1342 dvdd.n13 dvdd.n8 3.5845
R1343 dvdd.n13 dvdd.n12 3.1005
R1344 dvdd.n39 dvdd.n38 2.3255
R1345 dvdd.n40 dvdd.n1 0.317167
R1346 dvdd.n43 dvdd.n0 0.227778
R1347 dvdd.n44 dvdd 0.184693
R1348 dvdd.n42 dvdd.n1 0.153726
R1349 dvdd.n43 dvdd.n42 0.130913
R1350 dvdd.n38 dvdd.n37 0.129793
R1351 dvdd dvdd.n44 0.0827019
R1352 dvdd.n44 dvdd.n43 0.0726665
R1353 dvdd.n40 dvdd.n39 0.038
R1354 dvdd.n12 dvdd.n0 0.0212851
R1355 dvdd.n42 dvdd.n41 0.00788189
R1356 dvdd dvdd.n40 0.004875
R1357 dvdd.n41 dvdd 0.001125
R1358 dvdd.n41 dvdd 0.000992126
R1359 a_2982_4700.t1 a_2982_4700.n0 661.462
R1360 a_2982_4700.n0 a_2982_4700.t0 235.724
R1361 a_2982_4700.n0 a_2982_4700.t3 128.278
R1362 a_2982_4700.n0 a_2982_4700.t2 107.805
R1363 a_2982_4700.n1 a_2982_4700.t4 107.362
R1364 a_2982_4700.n1 a_2982_4700.t5 105.01
R1365 a_2982_4700.n0 a_2982_4700.n1 13.2005
R1366 dvss.n32 dvss.n16 2126.44
R1367 dvss.n37 dvss.n16 2126.44
R1368 dvss.n32 dvss.n17 2126.44
R1369 dvss.n37 dvss.n17 2126.44
R1370 dvss.n33 dvss.n28 1877.44
R1371 dvss.n27 dvss.n18 1836.74
R1372 dvss.n23 dvss.n19 1836.74
R1373 dvss.n27 dvss.n19 1836.74
R1374 dvss.n52 dvss.n11 1790.38
R1375 dvss.n51 dvss.n11 1790.38
R1376 dvss.n52 dvss.n12 1790.38
R1377 dvss.n51 dvss.n12 1790.38
R1378 dvss.n36 dvss.n35 1449.84
R1379 dvss.n48 dvss.n41 1407.97
R1380 dvss.n48 dvss.n47 1407.97
R1381 dvss.n42 dvss.n41 1407.97
R1382 dvss.n47 dvss.n42 1407.97
R1383 dvss.n28 dvss.t0 746.725
R1384 dvss.n34 dvss.n14 592.715
R1385 dvss.t5 dvss.n33 569.837
R1386 dvss.n23 dvss.n22 563.245
R1387 dvss.n46 dvss.t4 468.853
R1388 dvss.t2 dvss.n13 367.87
R1389 dvss.n34 dvss.t5 317.377
R1390 dvss.n30 dvss.n16 294.214
R1391 dvss.n47 dvss.n45 292.613
R1392 dvss.n25 dvss.n19 292.5
R1393 dvss.n19 dvss.t0 292.5
R1394 dvss.n21 dvss.n18 292.5
R1395 dvss.n47 dvss.n46 292.5
R1396 dvss.n44 dvss.n42 292.5
R1397 dvss.n42 dvss.t4 292.5
R1398 dvss.n43 dvss.n41 292.5
R1399 dvss.n41 dvss.n13 292.5
R1400 dvss.n49 dvss.n48 292.5
R1401 dvss.n48 dvss.t4 292.5
R1402 dvss.n51 dvss.n50 292.5
R1403 dvss.t2 dvss.n51 292.5
R1404 dvss.n53 dvss.n52 292.5
R1405 dvss.n52 dvss.t2 292.5
R1406 dvss.n17 dvss.n15 292.5
R1407 dvss.t5 dvss.n17 292.5
R1408 dvss.t5 dvss.n16 292.5
R1409 dvss.n36 dvss.n34 252.459
R1410 dvss.n55 dvss.t3 239.136
R1411 dvss.n1 dvss.t1 229.279
R1412 dvss.n35 dvss.n13 201.968
R1413 dvss.n27 dvss.n26 195
R1414 dvss.n28 dvss.n27 195
R1415 dvss.n24 dvss.n23 195
R1416 dvss.n12 dvss.n10 195
R1417 dvss.n46 dvss.n12 195
R1418 dvss.n11 dvss.n9 195
R1419 dvss.n35 dvss.n11 195
R1420 dvss.n22 dvss.n18 174.945
R1421 dvss.n38 dvss.n37 146.25
R1422 dvss.n37 dvss.n36 146.25
R1423 dvss.n32 dvss.n31 146.25
R1424 dvss.n33 dvss.n32 146.25
R1425 dvss.n31 dvss.n15 138.166
R1426 dvss.n53 dvss.n10 116.504
R1427 dvss.t2 dvss.t4 100.984
R1428 dvss.n22 dvss.t0 89.6975
R1429 dvss.n31 dvss.n30 86.5887
R1430 dvss.n25 dvss.n24 86.1306
R1431 dvss.n3 dvss.t6 84.1047
R1432 dvss.n24 dvss.n21 74.9169
R1433 dvss.n38 dvss.n15 59.6884
R1434 dvss.n40 dvss.n10 57.0178
R1435 dvss.n54 dvss.n53 53.0829
R1436 dvss.n45 dvss.n40 42.7428
R1437 dvss.n26 dvss.n25 41.1625
R1438 dvss.n45 dvss.n44 37.2564
R1439 dvss.n50 dvss.n39 31.8699
R1440 dvss.n44 dvss.n43 29.0402
R1441 dvss.n43 dvss.n39 26.2862
R1442 dvss.n20 dvss.n8 17.1865
R1443 dvss.n55 dvss.n54 14.0183
R1444 dvss.n21 dvss.n8 13.3694
R1445 dvss.n39 dvss.n14 11.3033
R1446 dvss.n49 dvss.n40 6.79341
R1447 dvss.n5 dvss.n2 5.813
R1448 dvss.n30 dvss.n29 5.6005
R1449 dvss.n54 dvss.n9 4.75646
R1450 dvss.n20 dvss.n1 4.6505
R1451 dvss.n26 dvss.n20 2.95435
R1452 dvss.n3 dvss.n2 2.6255
R1453 dvss.n29 dvss.n0 2.3255
R1454 dvss.n29 dvss.n14 1.88621
R1455 dvss.n56 dvss.n8 1.8479
R1456 dvss.n56 dvss.n55 1.50536
R1457 dvss.n50 dvss.n49 1.46336
R1458 dvss.n4 dvss.n3 1.2505
R1459 dvss.n5 dvss 0.8755
R1460 dvss.n4 dvss 0.583833
R1461 dvss.n7 dvss.n2 0.438
R1462 dvss.n14 dvss.n9 0.26472
R1463 dvss.n56 dvss 0.1955
R1464 dvss.n57 dvss.n1 0.170822
R1465 dvss.n58 dvss.n57 0.148685
R1466 dvss.n57 dvss.n7 0.142313
R1467 dvss.n7 dvss.n6 0.0735994
R1468 dvss.n39 dvss.n38 0.0592156
R1469 dvss.n6 dvss.n5 0.0415305
R1470 dvss.n57 dvss.n56 0.0277177
R1471 dvss.n58 dvss.n0 0.0276947
R1472 dvss.n6 dvss.n0 0.0200611
R1473 dvss.n6 dvss 0.0107339
R1474 dvss dvss.n58 0.00755645
R1475 dvss.n5 dvss.n4 0.0019313
R1476 dvss.n4 dvss 0.000977099
R1477 rc_osc_level_shifter_0.out_h rc_osc_level_shifter_0.out_h.t1 660.24
R1478 rc_osc_level_shifter_0.out_h rc_osc_level_shifter_0.out_h.t0 235.251
R1479 rc_osc_level_shifter_0.out_h rc_osc_level_shifter_0.out_h.t3 116.338
R1480 rc_osc_level_shifter_0.out_h.n0 rc_osc_level_shifter_0.out_h.t2 110.648
R1481 rc_osc_level_shifter_0.out_h rc_osc_level_shifter_0.out_h.t5 106.773
R1482 rc_osc_level_shifter_0.out_h.n0 rc_osc_level_shifter_0.out_h.t6 106.382
R1483 rc_osc_level_shifter_0.out_h.n0 rc_osc_level_shifter_0.out_h.t4 104.746
R1484 rc_osc_level_shifter_0.out_h rc_osc_level_shifter_0.out_h.n0 19.5701
R1485 a_1414_4786.n0 a_1414_4786.t3 237.433
R1486 a_1414_4786.n0 a_1414_4786.t2 235.407
R1487 a_1414_4786.t1 a_1414_4786.n0 233.657
R1488 a_1414_4786.n0 a_1414_4786.t7 111.246
R1489 a_1414_4786.n0 a_1414_4786.t4 105.537
R1490 a_1414_4786.n0 a_1414_4786.t0 104.177
R1491 a_1414_4786.n0 a_1414_4786.t6 104.175
R1492 a_1414_4786.n0 a_1414_4786.t9 104.175
R1493 a_1414_4786.n0 a_1414_4786.t5 104.175
R1494 a_1414_4786.n0 a_1414_4786.t8 104.175
R1495 a_514_7168.t0 a_514_7168.t1 245.351
R1496 dout dout.t2 243.404
R1497 dout.n0 dout.t0 229.669
R1498 dout.n0 dout.t1 171.274
R1499 dout dout.n0 2.52767
C0 a_6602_4786# dout 0.970428f
C1 avss a_514_9068# 0.305392f
C2 avss a_1344_7168# 0.239502f
C3 a_5826_9068# a_5494_9068# 0.307869f
C4 rc_osc_level_shifter_0.out_h a_3082_4788# 0.115135f
C5 rc_osc_level_shifter_0.out_h a_2526_4188# 0.106807f
C6 a_3834_9068# avss 0.142763f
C7 avss a_8170_1218# 0.158768f
C8 a_1012_7168# a_1344_7168# 0.307869f
C9 a_8366_5327# rc_osc_level_shifter_0.outb_h 0.202516f
C10 ena a_8366_5327# 0.117123f
C11 avss a_700_3118# 0.725274f
C12 a_4996_7168# a_4664_7168# 0.307869f
C13 a_9664_3118# a_9996_3118# 0.307869f
C14 a_6510_1218# a_6842_1218# 0.307869f
C15 avss a_8336_3118# 0.214531f
C16 avss a_5148_4788# 0.804644f
C17 a_7486_9068# a_7154_9068# 0.307869f
C18 a_6344_3118# a_6012_3118# 0.307869f
C19 a_4750_4788# a_5148_4788# 0.162171f
C20 a_9498_1218# avss 0.158768f
C21 a_2858_1218# avss 0.158903f
C22 avss a_2526_1218# 0.158903f
C23 a_3622_5653# a_3082_4788# 0.11132f
C24 a_3668_7168# avdd 0.547747f
C25 a_7672_3118# avss 0.216245f
C26 a_4000_7168# avdd 0.384982f
C27 avdd a_7598_4659# 0.401456f
C28 a_3336_7168# a_3668_7168# 0.307869f
C29 a_6842_1218# a_7174_1218# 0.307869f
C30 avss a_7652_7168# 0.243852f
C31 avss a_6158_9068# 0.142763f
C32 rc_osc_level_shifter_0.inb_l dout 0.168211f
C33 a_5992_7168# a_5660_7168# 0.307869f
C34 a_8814_9068# avss 0.142763f
C35 a_9332_3118# avss 0.208599f
C36 a_2692_3118# a_3024_3118# 0.307869f
C37 avss a_3082_4788# 0.767796f
C38 a_2008_7168# a_2340_7168# 0.307869f
C39 avss a_2526_4188# 0.660979f
C40 a_5992_7168# avdd 0.206045f
C41 avss a_4996_7168# 0.209517f
C42 a_3638_4788# rc_osc_level_shifter_0.outb_h 0.115253f
C43 a_6822_9068# a_7154_9068# 0.307869f
C44 avss dvdd 1.32271f
C45 avdd dout 0.101194f
C46 avss a_6656_7168# 0.209517f
C47 a_5992_7168# a_6324_7168# 0.307869f
C48 a_4996_7168# a_5328_7168# 0.307869f
C49 a_4750_4788# a_5470_5653# 0.111356f
C50 avss a_4664_7168# 0.209517f
C51 avss rc_osc_level_shifter_0.out_h 2.19553f
C52 ena rc_osc_level_shifter_0.outb_h 0.461732f
C53 avss a_7838_1218# 0.158768f
C54 a_4518_1218# a_4186_1218# 0.307869f
C55 a_4750_4788# rc_osc_level_shifter_0.out_h 0.155226f
C56 avss a_2174_9068# 0.142763f
C57 avss a_1530_1218# 0.158768f
C58 a_3638_4788# a_4194_4788# 0.365446f
C59 avss a_4684_3118# 0.256408f
C60 a_8004_3118# a_8336_3118# 0.307869f
C61 a_9312_7168# a_8980_7168# 0.307869f
C62 a_9478_9068# a_9146_9068# 0.307869f
C63 a_10681_5200# dout 0.224263f
C64 avss a_1178_9068# 0.142763f
C65 avss a_3356_3118# 0.63809f
C66 a_4036_4788# a_3638_4788# 0.162238f
C67 avss a_1364_3118# 0.280948f
C68 a_9332_3118# a_9664_3118# 0.307869f
C69 a_6988_7168# a_7320_7168# 0.307869f
C70 rc_osc_level_shifter_0.outb_h a_4194_4788# 0.124069f
C71 a_7672_3118# a_8004_3118# 0.307869f
C72 a_8316_7168# a_8648_7168# 0.307869f
C73 avss a_6676_3118# 0.723199f
C74 a_5182_1218# a_4850_1218# 0.307869f
C75 a_6178_1218# a_5846_1218# 0.307869f
C76 a_8814_9068# a_8482_9068# 0.307869f
C77 avss a_9976_7168# 0.144827f
C78 a_3190_1218# a_2858_1218# 0.307869f
C79 avss a_3854_1218# 0.158768f
C80 a_9166_1218# a_9498_1218# 0.307869f
C81 avss a_2672_7168# 0.209517f
C82 a_5680_3118# a_5348_3118# 0.307869f
C83 a_8668_3118# a_8336_3118# 0.307869f
C84 a_8648_7168# a_8980_7168# 0.307869f
C85 avss a_4750_4788# 0.857461f
C86 a_1012_7168# avss 0.239502f
C87 a_4830_9068# avss 0.142763f
C88 avss a_5328_7168# 0.209517f
C89 a_1510_9068# a_1842_9068# 0.307869f
C90 a_7598_4659# rc_osc_level_shifter_0.out_h 0.329503f
C91 a_2692_3118# a_2360_3118# 0.307869f
C92 a_1530_1218# a_1198_1218# 0.307869f
C93 avdd a_8366_5327# 0.528099f
C94 dvdd dout 0.536524f
C95 a_6602_4786# rc_osc_level_shifter_0.outb_h 0.183568f
C96 ena a_6602_4786# 0.523617f
C97 a_6490_9068# a_6158_9068# 0.307869f
C98 a_2028_3118# a_2360_3118# 0.307869f
C99 avss a_6444_4786# 0.405366f
C100 avss a_5514_1218# 0.158903f
C101 a_9332_3118# a_9000_3118# 0.307869f
C102 a_4518_1218# a_4850_1218# 0.307869f
C103 a_9644_7168# avdd 0.420324f
C104 a_1530_1218# a_1862_1218# 0.307869f
C105 a_9312_7168# avdd 0.206188f
C106 a_8814_9068# a_9146_9068# 0.307869f
C107 a_6012_3118# avss 0.539589f
C108 avss a_9664_3118# 0.208599f
C109 a_3668_7168# avss 0.209517f
C110 a_534_1218# a_866_1218# 0.307869f
C111 avss a_1198_1218# 0.158768f
C112 a_4000_7168# avss 0.209517f
C113 a_8502_1218# a_8834_1218# 0.307869f
C114 a_3480_4788# a_3082_4788# 0.161788f
C115 a_7838_1218# a_7506_1218# 0.307869f
C116 a_3834_9068# a_4166_9068# 0.307869f
C117 a_3638_4788# a_4238_5653# 0.111527f
C118 avss a_8150_9068# 0.142763f
C119 a_4592_4788# a_4194_4788# 0.161362f
C120 a_3004_7168# avdd 0.55108f
C121 rc_osc_level_shifter_0.inb_l rc_osc_level_shifter_0.outb_h 0.228327f
C122 ena rc_osc_level_shifter_0.inb_l 1.50031f
C123 a_3638_4788# avdd 0.824985f
C124 a_8482_9068# avss 0.142763f
C125 a_3004_7168# a_3336_7168# 0.307869f
C126 avss a_8004_3118# 0.215027f
C127 avss a_5992_7168# 0.209517f
C128 a_8648_7168# avdd 0.158636f
C129 avss a_1862_1218# 0.158903f
C130 a_10162_1218# a_9830_1218# 0.307869f
C131 avss a_680_7168# 0.238959f
C132 a_1676_7168# a_1344_7168# 0.307869f
C133 avss a_4498_9068# 0.142763f
C134 avdd rc_osc_level_shifter_0.outb_h 1.61593f
C135 ena avdd 1.61962f
C136 a_1012_7168# a_680_7168# 0.307869f
C137 a_10308_7168# a_9996_3118# 0.332125f
C138 a_4830_9068# a_4498_9068# 0.307869f
C139 a_3190_1218# avss 0.158903f
C140 a_10308_7168# rc_osc_level_shifter_0.inb_l 0.168314f
C141 a_4664_7168# a_4332_7168# 0.307869f
C142 a_3854_1218# a_4186_1218# 0.307869f
C143 a_9166_1218# avss 0.158768f
C144 avss a_4186_1218# 0.158768f
C145 a_6490_9068# avss 0.142763f
C146 avss a_7506_1218# 0.158768f
C147 avss a_2008_7168# 0.209517f
C148 avss a_9000_3118# 0.208599f
C149 a_8316_7168# a_7984_7168# 0.307869f
C150 a_4000_7168# a_3668_7168# 0.307869f
C151 a_6676_3118# a_7008_3118# 0.307869f
C152 avss a_8668_3118# 0.208599f
C153 a_8366_5327# rc_osc_level_shifter_0.out_h 0.102675f
C154 a_2028_3118# a_1696_3118# 0.307869f
C155 a_10308_7168# avdd 1.5149f
C156 avdd a_4194_4788# 0.827473f
C157 avss a_7008_3118# 0.337662f
C158 a_9810_9068# a_10142_9068# 0.307869f
C159 avss a_9146_9068# 0.142763f
C160 a_5826_9068# a_6158_9068# 0.307869f
C161 a_7818_9068# avss 0.142763f
C162 a_6988_7168# a_6656_7168# 0.307869f
C163 avss a_3480_4788# 0.752476f
C164 avss a_5680_3118# 0.677534f
C165 a_7672_3118# a_7340_3118# 0.307869f
C166 avss a_2924_4788# 0.817349f
C167 a_8482_9068# a_8150_9068# 0.307869f
C168 rc_osc_level_shifter_0.inb_l a_6602_4786# 0.903569f
C169 a_2526_1218# a_2194_1218# 0.307869f
C170 a_3522_1218# a_3854_1218# 0.307869f
C171 a_3638_4788# a_3082_4788# 0.378469f
C172 a_3522_1218# avss 0.158768f
C173 a_5162_9068# avss 0.142763f
C174 a_3502_9068# a_3170_9068# 0.307869f
C175 avss a_4332_7168# 0.209517f
C176 a_3170_9068# avdd 0.377892f
C177 a_5348_3118# a_5016_3118# 0.307869f
C178 a_5162_9068# a_4830_9068# 0.307869f
C179 a_8980_7168# avdd 0.198919f
C180 a_6602_4786# avdd 0.578691f
C181 rc_osc_level_shifter_0.outb_h a_3082_4788# 0.105461f
C182 a_4854_5653# a_4194_4788# 0.112519f
C183 a_3688_3118# a_4020_3118# 0.307869f
C184 a_3638_4788# rc_osc_level_shifter_0.out_h 0.131453f
C185 a_3024_3118# a_3356_3118# 0.307869f
C186 dvdd ena 1.36511f
C187 avss a_4850_1218# 0.158768f
C188 a_2506_9068# avdd 0.377892f
C189 a_4352_3118# a_4020_3118# 0.307869f
C190 a_9644_7168# a_9976_7168# 0.307869f
C191 a_6510_1218# avss 0.158903f
C192 a_6178_1218# avss 0.158892f
C193 a_4166_9068# avss 0.142763f
C194 a_9644_7168# avss 0.144844f
C195 a_6012_3118# a_5680_3118# 0.307869f
C196 a_5494_9068# avss 0.142763f
C197 a_9312_7168# avss 0.144844f
C198 rc_osc_level_shifter_0.out_h rc_osc_level_shifter_0.outb_h 3.38349f
C199 ena rc_osc_level_shifter_0.out_h 0.355894f
C200 a_6988_7168# avss 0.217519f
C201 a_9810_9068# a_9478_9068# 0.307869f
C202 a_7818_9068# a_8150_9068# 0.307869f
C203 avdd a_2340_7168# 0.399256f
C204 avss a_7154_9068# 0.142763f
C205 avss a_8834_1218# 0.158768f
C206 a_10308_7168# dvdd 0.994996f
C207 avss a_3024_3118# 0.739288f
C208 avss a_7174_1218# 0.158768f
C209 a_4000_7168# a_4332_7168# 0.307869f
C210 a_1510_9068# a_1178_9068# 0.307869f
C211 rc_osc_level_shifter_0.inb_l avdd 0.381808f
C212 a_5826_9068# avss 0.142763f
C213 a_3004_7168# avss 0.209517f
C214 avss a_1676_7168# 0.228829f
C215 a_9498_1218# a_9830_1218# 0.307869f
C216 rc_osc_level_shifter_0.out_h a_4194_4788# 0.145295f
C217 a_3004_7168# a_2672_7168# 0.307869f
C218 a_5660_7168# avdd 0.543399f
C219 avss a_7486_9068# 0.142763f
C220 avss a_3638_4788# 0.805426f
C221 avdd a_4238_5653# 0.701946f
C222 a_8668_3118# a_9000_3118# 0.307869f
C223 a_8648_7168# avss 0.148144f
C224 a_7320_7168# a_7652_7168# 0.307869f
C225 avss a_7340_3118# 0.220881f
C226 avss a_6842_1218# 0.158846f
C227 avss a_1510_9068# 0.142763f
C228 a_3336_7168# avdd 0.547747f
C229 avss rc_osc_level_shifter_0.outb_h 2.37072f
C230 avss ena 1.12459f
C231 avss a_2194_1218# 0.158903f
C232 a_3190_1218# a_3522_1218# 0.307869f
C233 dvdd a_6602_4786# 1.21653f
C234 a_4750_4788# rc_osc_level_shifter_0.outb_h 0.1288f
C235 a_700_3118# a_1032_3118# 0.307869f
C236 a_2692_3118# avss 0.739288f
C237 a_4684_3118# a_5016_3118# 0.307869f
C238 a_514_9068# a_846_9068# 0.307869f
C239 a_3834_9068# a_3502_9068# 0.307869f
C240 a_2028_3118# avss 0.739288f
C241 a_1842_9068# a_2174_9068# 0.307869f
C242 avdd a_700_3118# 0.308767f
C243 a_6602_4786# rc_osc_level_shifter_0.out_h 0.144369f
C244 a_8502_1218# a_8170_1218# 0.307869f
C245 a_10308_7168# a_9976_7168# 0.316348f
C246 a_7984_7168# a_7652_7168# 0.307869f
C247 ena a_6444_4786# 0.161553f
C248 a_6822_9068# avss 0.142763f
C249 avss a_4194_4788# 0.82682f
C250 a_10308_7168# avss 0.749668f
C251 avss a_534_1218# 0.322617f
C252 a_4750_4788# a_4194_4788# 0.385875f
C253 a_4166_9068# a_4498_9068# 0.307869f
C254 avdd a_4854_5653# 0.680997f
C255 avss a_4036_4788# 0.748363f
C256 a_2506_9068# a_2174_9068# 0.307869f
C257 a_8316_7168# avss 0.243852f
C258 avss a_5016_3118# 0.282044f
C259 a_10162_1218# avss 0.332866f
C260 dvdd rc_osc_level_shifter_0.inb_l 1.53482f
C261 avss a_2360_3118# 0.739288f
C262 a_7598_4659# rc_osc_level_shifter_0.outb_h 0.229013f
C263 a_3170_9068# avss 0.142763f
C264 avss a_1842_9068# 0.142763f
C265 a_9166_1218# a_8834_1218# 0.307869f
C266 avdd a_3082_4788# 0.817798f
C267 avss a_10142_9068# 0.304184f
C268 avss a_8980_7168# 0.144844f
C269 avss a_6602_4786# 0.609934f
C270 rc_osc_level_shifter_0.inb_l rc_osc_level_shifter_0.out_h 0.255748f
C271 avss a_866_1218# 0.158903f
C272 a_7320_7168# avss 0.243852f
C273 a_7174_1218# a_7506_1218# 0.307869f
C274 dvdd avdd 1.5343f
C275 avss a_9830_1218# 0.158768f
C276 a_2194_1218# a_1862_1218# 0.307869f
C277 avdd a_5470_5653# 0.763917f
C278 a_2008_7168# a_1676_7168# 0.307869f
C279 a_2858_1218# a_2526_1218# 0.307869f
C280 avss a_2506_9068# 0.142763f
C281 avss a_4592_4788# 0.748501f
C282 avss a_4020_3118# 0.255755f
C283 a_6324_7168# a_6656_7168# 0.307869f
C284 avdd rc_osc_level_shifter_0.out_h 2.36468f
C285 a_5162_9068# a_5494_9068# 0.307869f
C286 avss a_5846_1218# 0.158787f
C287 a_1032_3118# a_1364_3118# 0.307869f
C288 avss a_5182_1218# 0.158782f
C289 a_3688_3118# a_3356_3118# 0.307869f
C290 avss a_2340_7168# 0.209517f
C291 a_4684_3118# a_4352_3118# 0.307869f
C292 a_2672_7168# a_2340_7168# 0.307869f
C293 dvdd a_10681_5200# 0.244559f
C294 a_7818_9068# a_7486_9068# 0.307869f
C295 a_9810_9068# avss 0.142763f
C296 avss a_7984_7168# 0.243852f
C297 a_1178_9068# a_846_9068# 0.307869f
C298 avss a_9996_3118# 0.207783f
C299 a_7340_3118# a_7008_3118# 0.307869f
C300 a_7838_1218# a_8170_1218# 0.307869f
C301 a_3006_5653# avdd 0.816596f
C302 avss rc_osc_level_shifter_0.inb_l 0.882232f
C303 a_6344_3118# a_6676_3118# 0.307869f
C304 a_3622_5653# avdd 0.790633f
C305 a_1696_3118# a_1364_3118# 0.307869f
C306 a_5846_1218# a_5514_1218# 0.307869f
C307 avss a_1032_3118# 0.613897f
C308 a_1198_1218# a_866_1218# 0.307869f
C309 a_6510_1218# a_6178_1218# 0.307869f
C310 avss a_5660_7168# 0.209517f
C311 a_5514_1218# a_5182_1218# 0.307869f
C312 a_9478_9068# avss 0.142763f
C313 a_3688_3118# avss 0.272498f
C314 a_6344_3118# avss 0.739171f
C315 a_6822_9068# a_6490_9068# 0.307869f
C316 a_9312_7168# a_9644_7168# 0.307869f
C317 a_9976_7168# avdd 0.526222f
C318 a_5660_7168# a_5328_7168# 0.307869f
C319 a_3502_9068# avss 0.142763f
C320 avss a_4518_1218# 0.158768f
C321 avss avdd 0.256591p
C322 avss a_4352_3118# 0.254161f
C323 a_2672_7168# avdd 0.55108f
C324 avss a_846_9068# 0.142763f
C325 avdd a_4750_4788# 0.827529f
C326 a_8502_1218# avss 0.158768f
C327 a_3336_7168# avss 0.209517f
C328 avdd a_5328_7168# 0.435522f
C329 avss a_6324_7168# 0.209517f
C330 a_1696_3118# avss 0.530794f
C331 avss a_5348_3118# 0.669471f
C332 dout dvss 1.48439f
C333 ena dvss 1.28355f
C334 dvdd dvss 5.67086f
C335 avss dvss 7.015866f
C336 avdd dvss 0.302188p
C337 a_10162_1218# dvss 0.288134f
C338 a_9996_3118# dvss 0.233958f
C339 a_9830_1218# dvss 0.253248f
C340 a_9664_3118# dvss 0.233958f
C341 a_9498_1218# dvss 0.253248f
C342 a_9332_3118# dvss 0.233958f
C343 a_9166_1218# dvss 0.253248f
C344 a_9000_3118# dvss 0.233958f
C345 a_8834_1218# dvss 0.253248f
C346 a_8668_3118# dvss 0.233958f
C347 a_8502_1218# dvss 0.253248f
C348 a_8336_3118# dvss 0.233958f
C349 a_8170_1218# dvss 0.253248f
C350 a_8004_3118# dvss 0.233958f
C351 a_7838_1218# dvss 0.253248f
C352 a_7672_3118# dvss 0.233958f
C353 a_7506_1218# dvss 0.253248f
C354 a_7340_3118# dvss 0.233958f
C355 a_7174_1218# dvss 0.253248f
C356 a_7008_3118# dvss 0.233958f
C357 a_6842_1218# dvss 0.253248f
C358 a_6676_3118# dvss 0.233958f
C359 a_6510_1218# dvss 0.253248f
C360 a_6344_3118# dvss 0.233958f
C361 a_6178_1218# dvss 0.253248f
C362 a_6012_3118# dvss 0.233958f
C363 a_5846_1218# dvss 0.253248f
C364 a_5680_3118# dvss 0.233958f
C365 a_5514_1218# dvss 0.253248f
C366 a_5348_3118# dvss 0.233958f
C367 a_5182_1218# dvss 0.253248f
C368 a_5016_3118# dvss 0.233958f
C369 a_4850_1218# dvss 0.253248f
C370 a_4684_3118# dvss 0.233958f
C371 a_4518_1218# dvss 0.253248f
C372 a_4352_3118# dvss 0.233958f
C373 a_4186_1218# dvss 0.253248f
C374 a_4020_3118# dvss 0.233958f
C375 a_3854_1218# dvss 0.253248f
C376 a_3688_3118# dvss 0.233958f
C377 a_3522_1218# dvss 0.253248f
C378 a_3356_3118# dvss 0.233958f
C379 a_3190_1218# dvss 0.253248f
C380 a_3024_3118# dvss 0.233958f
C381 a_2858_1218# dvss 0.253248f
C382 a_2692_3118# dvss 0.233958f
C383 a_2526_1218# dvss 0.253248f
C384 a_2360_3118# dvss 0.233958f
C385 a_2194_1218# dvss 0.253248f
C386 a_2028_3118# dvss 0.233958f
C387 a_1862_1218# dvss 0.253248f
C388 a_1696_3118# dvss 0.233958f
C389 a_1530_1218# dvss 0.253248f
C390 a_1364_3118# dvss 0.233958f
C391 a_1198_1218# dvss 0.253248f
C392 a_1032_3118# dvss 0.236415f
C393 a_866_1218# dvss 0.253248f
C394 a_700_3118# dvss 0.241208f
C395 a_534_1218# dvss 0.288266f
C396 rc_osc_level_shifter_0.outb_h dvss 3.514437f
C397 rc_osc_level_shifter_0.inb_l dvss 1.19529f
C398 a_6602_4786# dvss 0.840191f
C399 a_4750_4788# dvss 0.148139f
C400 a_4194_4788# dvss 0.146283f
C401 a_3638_4788# dvss 0.145977f
C402 a_3082_4788# dvss 0.145888f
C403 rc_osc_level_shifter_0.out_h dvss 4.252511f
C404 a_10308_7168# dvss 2.36722f
C405 a_10142_9068# dvss 0.289538f
C406 a_9976_7168# dvss 0.233244f
C407 a_9810_9068# dvss 0.25332f
C408 a_9644_7168# dvss 0.232864f
C409 a_9478_9068# dvss 0.25332f
C410 a_9312_7168# dvss 0.232864f
C411 a_9146_9068# dvss 0.25332f
C412 a_8980_7168# dvss 0.232864f
C413 a_8814_9068# dvss 0.25332f
C414 a_8648_7168# dvss 0.234983f
C415 a_8482_9068# dvss 0.25332f
C416 a_8316_7168# dvss 0.232864f
C417 a_8150_9068# dvss 0.25332f
C418 a_7984_7168# dvss 0.232864f
C419 a_7818_9068# dvss 0.25332f
C420 a_7652_7168# dvss 0.232864f
C421 a_7486_9068# dvss 0.25332f
C422 a_7320_7168# dvss 0.232864f
C423 a_7154_9068# dvss 0.25332f
C424 a_6988_7168# dvss 0.232864f
C425 a_6822_9068# dvss 0.25332f
C426 a_6656_7168# dvss 0.232864f
C427 a_6490_9068# dvss 0.25332f
C428 a_6324_7168# dvss 0.232864f
C429 a_6158_9068# dvss 0.25332f
C430 a_5992_7168# dvss 0.232864f
C431 a_5826_9068# dvss 0.25332f
C432 a_5660_7168# dvss 0.232864f
C433 a_5494_9068# dvss 0.25332f
C434 a_5328_7168# dvss 0.232864f
C435 a_5162_9068# dvss 0.25332f
C436 a_4996_7168# dvss 0.232864f
C437 a_4830_9068# dvss 0.25332f
C438 a_4664_7168# dvss 0.232864f
C439 a_4498_9068# dvss 0.25332f
C440 a_4332_7168# dvss 0.232864f
C441 a_4166_9068# dvss 0.25332f
C442 a_4000_7168# dvss 0.232864f
C443 a_3834_9068# dvss 0.25332f
C444 a_3668_7168# dvss 0.232864f
C445 a_3502_9068# dvss 0.25332f
C446 a_3336_7168# dvss 0.232864f
C447 a_3170_9068# dvss 0.25332f
C448 a_3004_7168# dvss 0.232864f
C449 a_2672_7168# dvss 0.232864f
C450 a_2506_9068# dvss 0.25332f
C451 a_2340_7168# dvss 0.232864f
C452 a_2174_9068# dvss 0.25332f
C453 a_2008_7168# dvss 0.232864f
C454 a_1842_9068# dvss 0.25332f
C455 a_1676_7168# dvss 0.232864f
C456 a_1510_9068# dvss 0.25332f
C457 a_1344_7168# dvss 0.232864f
C458 a_1178_9068# dvss 0.25332f
C459 a_1012_7168# dvss 0.232864f
C460 a_846_9068# dvss 0.25332f
C461 a_680_7168# dvss 0.232864f
C462 a_514_9068# dvss 0.289263f
C463 a_514_7168.t0 dvss 2.0228f
C464 a_1414_4786.n0 dvss 5.92504f
C465 a_1414_4786.t4 dvss 0.343122f
C466 a_1414_4786.t6 dvss 0.337945f
C467 a_1414_4786.t9 dvss 0.337945f
C468 a_1414_4786.t5 dvss 0.337945f
C469 a_1414_4786.t8 dvss 0.337945f
C470 a_1414_4786.t7 dvss 0.337945f
C471 a_1414_4786.t0 dvss 0.337946f
C472 rc_osc_level_shifter_0.out_h.n0 dvss 3.00052f
C473 rc_osc_level_shifter_0.out_h.t5 dvss 0.221005f
C474 rc_osc_level_shifter_0.out_h.t3 dvss 0.257597f
C475 rc_osc_level_shifter_0.out_h.t6 dvss 0.21472f
C476 rc_osc_level_shifter_0.out_h.t4 dvss 0.209426f
C477 rc_osc_level_shifter_0.out_h.t2 dvss 0.235108f
C478 a_2982_4700.n0 dvss 1.53467f
C479 a_2982_4700.t2 dvss 0.117719f
C480 a_2982_4700.t3 dvss 0.174566f
C481 a_2982_4700.t4 dvss 0.116691f
C482 a_2982_4700.t5 dvss 0.110026f
C483 a_2982_4700.n1 dvss 0.702349f
C484 rc_osc_level_shifter_0.outb_h.n0 dvss 1.70946f
C485 rc_osc_level_shifter_0.outb_h.t2 dvss 0.427686f
C486 rc_osc_level_shifter_0.outb_h.t3 dvss 0.236427f
C487 rc_osc_level_shifter_0.outb_h.t4 dvss 0.204773f
C488 avdd.n0 dvss -2.08361f
C489 avdd.n1 dvss 0.121888f
C490 avdd.n2 dvss 0.231852f
C491 avdd.n3 dvss 0.115726f
C492 avdd.n4 dvss 0.115726f
C493 avdd.n5 dvss 1.36105f
C494 avdd.n6 dvss 0.115795f
C495 avdd.n7 dvss 0.115795f
C496 avdd.n8 dvss 1.38162f
C497 avdd.n9 dvss 0.55782f
C498 avdd.n10 dvss 0.176696f
C499 avdd.n11 dvss 0.115795f
C500 avdd.n12 dvss 0.115795f
C501 avdd.t26 dvss 0.730238f
C502 avdd.n13 dvss 0.115795f
C503 avdd.n14 dvss 0.115726f
C504 avdd.n15 dvss 0.129196f
C505 avdd.n16 dvss 0.973651f
C506 avdd.n17 dvss 1.25683f
C507 avdd.n18 dvss 0.768135f
C508 avdd.n19 dvss 0.689468f
C509 avdd.n20 dvss 0.793282f
C510 avdd.n21 dvss 0.79312f
C511 avdd.n22 dvss 3.21735f
C512 avdd.n23 dvss 11.5836f
C513 avdd.n24 dvss 2.70915f
C514 avdd.n25 dvss 4.64888f
C515 avdd.n26 dvss 2.70898f
C516 avdd.n27 dvss 5.13893f
C517 avdd.n28 dvss 0.897805f
C518 avdd.n29 dvss 0.905036f
C519 avdd.n30 dvss 2.93578f
C520 avdd.n31 dvss 1.66127f
C521 avdd.n32 dvss 1.10425f
C522 avdd.n33 dvss 3.29474f
C523 avdd.n34 dvss 0.685206f
C524 avdd.n35 dvss 0.431773f
C525 avdd.n36 dvss 0.431773f
C526 avdd.n37 dvss 0.224995f
C527 avdd.n41 dvss 0.2455f
C528 avdd.n42 dvss 0.115726f
C529 avdd.n44 dvss 1.1933f
C530 avdd.n45 dvss 0.115726f
C531 avdd.n47 dvss 1.2614f
C532 avdd.n49 dvss 0.156254f
C533 avdd.n56 dvss 1.2614f
C534 avdd.n60 dvss 0.242434f
C535 avdd.n66 dvss 0.156699f
C536 avdd.n67 dvss 0.115726f
C537 avdd.n68 dvss 0.115726f
C538 avdd.n69 dvss 1.1933f
C539 avdd.n70 dvss 0.115795f
C540 avdd.n71 dvss 1.1933f
C541 avdd.n72 dvss 0.115795f
C542 avdd.n73 dvss 0.115726f
C543 avdd.n74 dvss 0.115726f
C544 avdd.n77 dvss 0.156254f
C545 avdd.n78 dvss 0.115726f
C546 avdd.n79 dvss 0.115726f
C547 avdd.n80 dvss 1.1933f
C548 avdd.n81 dvss 0.115795f
C549 avdd.n82 dvss 0.115795f
C550 avdd.n83 dvss 1.1933f
C551 avdd.n84 dvss 0.126714f
C552 avdd.n85 dvss 0.115726f
C553 avdd.n88 dvss 0.156699f
C554 avdd.n89 dvss 0.115726f
C555 avdd.n90 dvss 0.115726f
C556 avdd.n91 dvss 1.1933f
C557 avdd.n92 dvss 0.115795f
C558 avdd.n93 dvss 1.1933f
C559 avdd.n94 dvss 0.115795f
C560 avdd.n95 dvss 0.115726f
C561 avdd.n96 dvss 0.115726f
C562 avdd.n97 dvss 1.24126f
C563 avdd.n99 dvss 0.431773f
C564 avdd.n102 dvss 0.126714f
C565 avdd.n103 dvss 0.115795f
C566 avdd.n104 dvss 0.115726f
C567 avdd.n105 dvss 0.115726f
C568 avdd.n106 dvss 1.1933f
C569 avdd.n107 dvss 0.115795f
C570 avdd.n108 dvss 1.1933f
C571 avdd.n109 dvss 0.115726f
C572 avdd.n110 dvss 0.115726f
C573 avdd.n113 dvss 0.164237f
C574 avdd.n115 dvss 0.115726f
C575 avdd.n116 dvss 1.2614f
C576 avdd.n117 dvss 0.115795f
C577 avdd.n118 dvss 0.115795f
C578 avdd.n119 dvss 1.1933f
C579 avdd.n121 dvss 0.126714f
C580 avdd.n122 dvss 0.115726f
C581 avdd.n124 dvss 0.185829f
C582 avdd.n125 dvss 0.115726f
C583 avdd.n126 dvss 1.01564f
C584 avdd.n128 dvss 0.346841f
C585 avdd.n129 dvss 0.129485f
C586 avdd.n130 dvss 1.16261f
C587 avdd.n131 dvss 0.135804f
C588 avdd.n132 dvss 1.0189f
C589 avdd.n133 dvss 0.270881f
C590 avdd.n135 dvss 0.115726f
C591 avdd.n137 dvss 0.156699f
C592 avdd.n138 dvss 0.147904f
C593 avdd.n140 dvss 0.156699f
C594 avdd.n141 dvss 0.156699f
C595 avdd.n142 dvss 0.147904f
C596 avdd.n143 dvss 0.283775f
C597 avdd.n144 dvss 0.288007f
C598 avdd.n145 dvss 0.293831f
C599 avdd.n146 dvss 0.138272f
C600 avdd.t27 dvss 1.09994f
C601 avdd.n147 dvss 0.138272f
C602 avdd.n149 dvss 0.762362f
C603 avdd.n150 dvss 0.464273f
C604 avdd.n151 dvss 0.147904f
C605 avdd.t9 dvss 1.2614f
C606 avdd.n154 dvss 0.201791f
C607 avdd.n157 dvss 0.220764f
C608 avdd.n158 dvss 0.432679f
C609 avdd.n159 dvss 2.19906f
C610 avdd.n160 dvss 0.635524f
C611 avdd.n161 dvss 0.431773f
C612 avdd.n162 dvss 0.209347f
C613 avdd.n163 dvss 0.224995f
C614 avdd.n164 dvss 0.108537f
C615 avdd.t12 dvss 1.2614f
C616 avdd.n167 dvss 0.147904f
C617 avdd.n168 dvss 0.156254f
C618 avdd.n169 dvss 0.156254f
C619 avdd.n170 dvss 0.109035f
C620 avdd.n171 dvss 0.156254f
C621 avdd.n172 dvss 0.147904f
C622 avdd.n173 dvss 0.115795f
C623 avdd.t0 dvss 1.2614f
C624 avdd.n174 dvss 0.115795f
C625 avdd.n175 dvss 0.108537f
C626 avdd.n176 dvss 0.224995f
C627 avdd.n177 dvss 0.209347f
C628 avdd.n179 dvss 0.126714f
C629 avdd.n180 dvss 0.108537f
C630 avdd.n182 dvss 0.209347f
C631 avdd.n183 dvss 0.224995f
C632 avdd.n185 dvss 0.156254f
C633 avdd.n186 dvss 0.121171f
C634 avdd.n187 dvss 0.115795f
C635 avdd.t1 dvss 1.2614f
C636 avdd.n188 dvss 0.115795f
C637 avdd.n189 dvss 0.147904f
C638 avdd.n190 dvss 0.156699f
C639 avdd.n191 dvss 0.156699f
C640 avdd.n192 dvss 0.147904f
C641 avdd.n193 dvss 0.156699f
C642 avdd.n194 dvss 0.115726f
C643 avdd.n196 dvss 0.108537f
C644 avdd.n198 dvss 0.126714f
C645 avdd.n199 dvss 0.209347f
C646 avdd.n200 dvss 0.224995f
C647 avdd.n201 dvss 0.108537f
C648 avdd.n202 dvss 0.115795f
C649 avdd.t3 dvss 1.2614f
C650 avdd.n203 dvss 0.115795f
C651 avdd.n204 dvss 0.147904f
C652 avdd.n205 dvss 0.156254f
C653 avdd.n206 dvss 0.156254f
C654 avdd.n208 dvss 0.156254f
C655 avdd.n209 dvss 0.147904f
C656 avdd.n210 dvss 0.115795f
C657 avdd.t5 dvss 1.2614f
C658 avdd.n211 dvss 0.115795f
C659 avdd.n212 dvss 0.147904f
C660 avdd.n213 dvss 0.156699f
C661 avdd.n214 dvss 0.156699f
C662 avdd.n215 dvss 0.147904f
C663 avdd.n216 dvss 0.164673f
C664 avdd.n217 dvss 0.146032f
C665 avdd.n218 dvss 0.162822f
C666 avdd.n220 dvss 0.115726f
C667 avdd.n221 dvss 0.268745f
C668 avdd.n223 dvss 1.1933f
C669 avdd.n225 dvss 0.115726f
C670 avdd.n226 dvss 0.276934f
C671 avdd.n227 dvss 0.367379f
C672 avdd.n228 dvss 0.252777f
C673 avdd.n229 dvss 0.123254f
C674 avdd.t17 dvss 1.2614f
C675 avdd.n235 dvss 0.229993f
C676 avdd.n236 dvss 0.209218f
C677 avdd.n237 dvss 0.184173f
C678 avdd.n238 dvss 0.503485f
C679 avdd.n239 dvss 0.10651f
C680 avdd.n240 dvss 0.122508f
C681 avdd.t7 dvss 1.2614f
C682 avdd.n244 dvss 0.171732f
C683 avdd.n245 dvss 0.147904f
C684 avdd.t14 dvss 1.2614f
C685 avdd.n248 dvss 0.108537f
C686 avdd.n249 dvss 0.126714f
C687 avdd.n250 dvss 0.209347f
C688 avdd.n251 dvss 0.580069f
C689 avdd.n252 dvss 1.1296f
C690 avdd.n253 dvss 1.615f
C691 avdd.n254 dvss 7.8968f
C692 avdd.t21 dvss 0.129222f
C693 avdd.n255 dvss 9.88555f
C694 avdd.n256 dvss 7.06723f
C695 avdd.n257 dvss 19.265501f
C696 avdd.n258 dvss 15.564799f
C697 avdd.n259 dvss 13.776f
C698 avdd.n260 dvss 2.25701f
C699 avdd.n261 dvss 0.677275f
C700 avdd.n262 dvss 1.80429f
C701 avdd.n263 dvss 1.52665f
C702 avdd.n264 dvss 6.53464f
C703 avdd.n265 dvss 11.5829f
C704 avdd.n266 dvss 13.779799f
C705 avdd.n267 dvss 3.19564f
C706 avdd.n268 dvss 2.77059f
C707 avdd.n269 dvss 3.83712f
C708 avdd.n270 dvss 2.10894f
C709 avdd.n271 dvss 1.52601f
C710 avdd.n272 dvss 6.532f
C711 avdd.n273 dvss 2.50428f
C712 avdd.n274 dvss 3.7174f
C713 avdd.n275 dvss 1.56692f
C714 avdd.n276 dvss 0.66748f
C715 avdd.n277 dvss 0.878617f
C716 avdd.n278 dvss 1.27507f
C717 avdd.n279 dvss 0.743135f
C718 avdd.n280 dvss 0.157445f
C719 avdd.n281 dvss 0.125229f
C720 avdd.n283 dvss 0.121499f
C721 avdd.n284 dvss 0.3041f
C722 avdd.n285 dvss 0.211577f
C723 avdd.n286 dvss 0.115726f
C724 avdd.n287 dvss 0.730238f
C725 avdd.t24 dvss 0.730238f
C726 avdd.n288 dvss 0.115795f
C727 avdd.n289 dvss 0.253916f
C728 avdd.n290 dvss 0.140383f
C729 avdd.n291 dvss 0.2387f
C730 avdd.n292 dvss 0.115726f
C731 avdd.n293 dvss 0.730238f
C732 avdd.n294 dvss 0.651386f
C733 avdd.n295 dvss 0.115726f
C734 avdd.n296 dvss 0.108537f
C735 avdd.n297 dvss 0.115726f
C736 avdd.n298 dvss 0.132815f
C737 avdd.n299 dvss 0.275722f
C738 avdd.n300 dvss 0.174423f
C739 avdd.n301 dvss 0.115726f
C740 avdd.n302 dvss 0.205075f
C741 avdd.n303 dvss 0.302734f
C742 avdd.n304 dvss 0.210837f
C743 avdd.n305 dvss 0.115795f
C744 avdd.t23 dvss 1.4551f
C745 avdd.n306 dvss 0.115795f
C746 avdd.n307 dvss 0.132308f
C747 avdd.n308 dvss 0.155396f
C748 a_1538_5653.n0 dvss 5.44118f
C749 a_1538_5653.n1 dvss 2.03869f
C750 a_1538_5653.t6 dvss 0.272024f
C751 a_1538_5653.t10 dvss 0.272094f
C752 a_1538_5653.t17 dvss 0.272094f
C753 a_1538_5653.t16 dvss 0.272094f
C754 a_1538_5653.t18 dvss 0.272094f
C755 a_1538_5653.t14 dvss 0.272094f
C756 a_1538_5653.t15 dvss 0.272094f
C757 a_1538_5653.t4 dvss 0.284083f
C758 a_1538_5653.t0 dvss 0.272024f
C759 a_1538_5653.t2 dvss 0.272019f
C760 a_1538_5653.t8 dvss 0.272019f
C761 avss.n0 dvss 2.58818f
C762 avss.n1 dvss 1.19805f
C763 avss.n2 dvss 1.73103f
C764 avss.n3 dvss 0.516994f
C765 avss.n4 dvss 0.516994f
C766 avss.t2 dvss 1.23687f
C767 avss.t123 dvss 0.781297f
C768 avss.n5 dvss 0.516994f
C769 avss.n6 dvss 0.516994f
C770 avss.n7 dvss 1.74084f
C771 avss.n8 dvss 1.42542f
C772 avss.n9 dvss 0.371052f
C773 avss.n10 dvss 0.314829f
C774 avss.n11 dvss 0.277174f
C775 avss.n12 dvss 1.42186f
C776 avss.t25 dvss 1.09552f
C777 avss.t125 dvss 1.09141f
C778 avss.t98 dvss 1.09141f
C779 avss.t41 dvss 1.09141f
C780 avss.t73 dvss 1.09141f
C781 avss.t77 dvss 1.09141f
C782 avss.t72 dvss 1.09141f
C783 avss.t63 dvss 1.09141f
C784 avss.t11 dvss 1.09141f
C785 avss.t56 dvss 1.09141f
C786 avss.t69 dvss 1.16047f
C787 avss.t117 dvss 1.15831f
C788 avss.t132 dvss 1.19495f
C789 avss.t129 dvss 1.19495f
C790 avss.t119 dvss 1.19495f
C791 avss.t32 dvss 0.925005f
C792 avss.t71 dvss 1.19535f
C793 avss.t19 dvss 1.19535f
C794 avss.t101 dvss 1.19535f
C795 avss.t130 dvss 1.19535f
C796 avss.t1 dvss 1.19535f
C797 avss.t54 dvss 1.19535f
C798 avss.t3 dvss 1.19535f
C799 avss.t17 dvss 1.19535f
C800 avss.t34 dvss 1.19535f
C801 avss.t49 dvss 1.19535f
C802 avss.t109 dvss 1.19535f
C803 avss.t42 dvss 1.19535f
C804 avss.t61 dvss 1.19535f
C805 avss.t22 dvss 1.19535f
C806 avss.t141 dvss 1.19535f
C807 avss.t66 dvss 1.19535f
C808 avss.t26 dvss 1.19535f
C809 avss.t35 dvss 1.19535f
C810 avss.t120 dvss 1.19535f
C811 avss.t78 dvss 1.19535f
C812 avss.t21 dvss 1.19535f
C813 avss.t58 dvss 1.19535f
C814 avss.t53 dvss 1.19535f
C815 avss.t43 dvss 1.19535f
C816 avss.t27 dvss 1.19535f
C817 avss.t14 dvss 1.19535f
C818 avss.t136 dvss 0.896512f
C819 avss.n13 dvss 0.597674f
C820 avss.t104 dvss 0.896512f
C821 avss.t80 dvss 1.19535f
C822 avss.t74 dvss 1.22921f
C823 avss.t45 dvss 1.16094f
C824 avss.t67 dvss 1.19495f
C825 avss.t13 dvss 1.19495f
C826 avss.t108 dvss 1.19495f
C827 avss.t15 dvss 1.19495f
C828 avss.t111 dvss 1.19495f
C829 avss.t116 dvss 1.19495f
C830 avss.t140 dvss 1.19495f
C831 avss.t40 dvss 1.19495f
C832 avss.t30 dvss 1.19495f
C833 avss.t16 dvss 0.867417f
C834 avss.n14 dvss 1.00806f
C835 avss.n19 dvss 0.158124f
C836 avss.n20 dvss 0.411624f
C837 avss.n22 dvss 0.929261f
C838 avss.n23 dvss 0.107625f
C839 avss.t121 dvss 1.25509f
C840 avss.t75 dvss 1.10469f
C841 avss.n27 dvss 0.136675f
C842 avss.n29 dvss 0.545869f
C843 avss.n33 dvss 0.448821f
C844 avss.n37 dvss 0.794165f
C845 avss.n41 dvss 0.315624f
C846 avss.n42 dvss 0.626832f
C847 avss.n43 dvss 0.381113f
C848 avss.n50 dvss 0.178853f
C849 avss.t112 dvss 1.11161f
C850 avss.t110 dvss 1.11161f
C851 avss.t124 dvss 1.11161f
C852 avss.t37 dvss 1.02811f
C853 avss.n66 dvss 0.178853f
C854 avss.n67 dvss 1.3941f
C855 avss.t105 dvss 1.11161f
C856 avss.t113 dvss 0.986362f
C857 avss.n81 dvss 0.165138f
C858 avss.t7 dvss 1.04899f
C859 avss.t64 dvss 1.30471f
C860 avss.n84 dvss 0.866328f
C861 avss.t128 dvss 1.11161f
C862 avss.n86 dvss 0.179651f
C863 avss.n87 dvss 0.240378f
C864 avss.n88 dvss 0.207163f
C865 avss.n89 dvss 0.141819f
C866 avss.n90 dvss 2.26925f
C867 avss.t86 dvss 0.965486f
C868 avss.t118 dvss 1.11161f
C869 avss.n98 dvss 0.866328f
C870 avss.t138 dvss 0.67845f
C871 avss.n99 dvss 0.866328f
C872 avss.t68 dvss 0.908079f
C873 avss.t24 dvss 1.09596f
C874 avss.t31 dvss 1.06986f
C875 avss.t96 dvss 0.866328f
C876 avss.n105 dvss 0.125574f
C877 avss.n106 dvss 0.133792f
C878 avss.n107 dvss 0.216153f
C879 avss.n108 dvss 0.216236f
C880 avss.t9 dvss 1.01246f
C881 avss.n113 dvss 0.824577f
C882 avss.n114 dvss 0.720201f
C883 avss.t6 dvss 0.866328f
C884 avss.n130 dvss 0.866328f
C885 avss.t126 dvss 0.67845f
C886 avss.n131 dvss 0.866328f
C887 avss.t10 dvss 1.00724f
C888 avss.t55 dvss 1.11161f
C889 avss.t133 dvss 0.94983f
C890 avss.n142 dvss 0.761951f
C891 avss.t134 dvss 0.970705f
C892 avss.n143 dvss 0.782827f
C893 avss.t29 dvss 1.11161f
C894 avss.n153 dvss 0.866328f
C895 avss.t106 dvss 0.67845f
C896 avss.n154 dvss 0.866328f
C897 avss.t107 dvss 0.99158f
C898 avss.t84 dvss 0.928954f
C899 avss.n166 dvss 0.741076f
C900 avss.n167 dvss 0.803702f
C901 avss.n170 dvss 0.304909f
C902 avss.n177 dvss 0.866328f
C903 avss.t70 dvss 0.67845f
C904 avss.n178 dvss 0.866328f
C905 avss.t82 dvss 1.11161f
C906 avss.t90 dvss 0.866328f
C907 avss.t88 dvss 0.866328f
C908 avss.n193 dvss 0.682246f
C909 avss.n194 dvss 2.41946f
C910 avss.n195 dvss 0.454528f
C911 avss.n196 dvss 0.648808f
C912 avss.n197 dvss 1.42629f
C913 avss.n198 dvss 0.604748f
C914 avss.n199 dvss 1.21333f
C915 avss.t65 dvss 1.58912f
C916 avss.t122 dvss 1.20636f
C917 avss.t8 dvss 1.24572f
C918 avss.t36 dvss 1.24572f
C919 avss.t18 dvss 1.24572f
C920 avss.t12 dvss 1.24572f
C921 avss.t93 dvss 1.24572f
C922 avss.t85 dvss 1.25583f
C923 avss.t137 dvss 1.10975f
C924 avss.t38 dvss 1.08981f
C925 avss.t60 dvss 1.08981f
C926 avss.t81 dvss 1.08981f
C927 avss.t5 dvss 1.08981f
C928 avss.t114 dvss 1.08981f
C929 avss.t131 dvss 1.08981f
C930 avss.t79 dvss 1.08981f
C931 avss.t62 dvss 1.08981f
C932 avss.t76 dvss 1.08981f
C933 avss.t135 dvss 1.08524f
C934 avss.n200 dvss 1.29791f
C935 avss.n201 dvss 0.897688f
C936 avss.n202 dvss 0.954135f
C937 avss.n203 dvss 5.57064f
C938 avss.n204 dvss 7.23255f
C939 avss.n205 dvss 4.63454f
C940 avss.n206 dvss 8.828441f
C941 avss.n207 dvss 2.96518f
C942 avss.n208 dvss 0.409181f
C943 avss.n209 dvss 1.44532f
C944 avss.n210 dvss 1.12451f
C945 avss.n211 dvss 4.53165f
C946 avss.n212 dvss 0.222922f
C947 avss.n213 dvss 0.136f
C948 avss.n214 dvss 0.11799f
C949 avss.t46 dvss 0.866328f
C950 avss.n218 dvss 0.150388f
C951 avss.t33 dvss 0.866328f
C952 avss.n228 dvss 0.178853f
C953 avss.n229 dvss 0.537382f
C954 avss.n230 dvss 0.178853f
C955 avss.t94 dvss 0.866328f
C956 avss.t50 dvss 0.866328f
C957 avss.n245 dvss 0.178853f
C958 avss.n246 dvss 0.404387f
C959 avss.n247 dvss 0.293471f
C960 avss.n248 dvss 0.178853f
C961 avss.n252 dvss 0.288229f
C962 avss.n254 dvss 0.433164f
C963 avss.t83 dvss 1.28384f
C964 avss.t39 dvss 1.73266f
C965 avss.t139 dvss 1.73266f
C966 avss.t28 dvss 1.73266f
C967 avss.t4 dvss 1.52282f
C968 avss.n256 dvss 0.860449f
C969 avss.t48 dvss 1.06838f
C970 avss.t127 dvss 0.897234f
C971 avss.t87 dvss 0.860929f
C972 avss.n259 dvss 0.100993f
C973 avss.n260 dvss 0.145906f
C974 avss.n261 dvss 0.137634f
C975 avss.n263 dvss 0.860931f
C976 avss.t44 dvss 1.4418f
C977 avss.t57 dvss 1.3277f
C978 avss.n264 dvss 1.58397f
C979 avss.t51 dvss 0.751312f
C980 avss.n266 dvss 1.16234f
C981 avss.n267 dvss 0.159237f
C982 avss.n268 dvss 0.108026f
C983 avss.n271 dvss 0.13778f
C984 avss.t102 dvss 0.853918f
C985 avss.n277 dvss 0.146277f
C986 avss.n280 dvss 0.174153f
C987 avss.n282 dvss 2.89458f
C988 avss.n283 dvss 0.104412f
C989 avss.n284 dvss 0.873843f
C990 avss.n285 dvss 1.79069f
C991 avss.n286 dvss 3.96852f
C992 avss.n287 dvss 1.54188f
C993 avss.t0 dvss 1.20907f
C994 avss.t20 dvss 1.01173f
C995 avss.n288 dvss 2.25665f
C996 avss.n289 dvss 2.5253f
C997 avss.t23 dvss 1.36212f
C998 avss.t59 dvss 1.81948f
C999 avss.n290 dvss 2.14362f
C1000 avss.n291 dvss 0.97592f
C1001 avss.n292 dvss 0.681449f
C1002 avss.n293 dvss 1.41609f
.ends

